module Gate();

wire a, b, z;

nand NAND2_X1 (z, a, b);

endmodule
