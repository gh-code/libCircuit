module empty();
wire a;
endmodule
