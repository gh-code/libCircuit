
module ethernet_syn_comb ( wb_dat_i_0, wb_dat_i_1, wb_dat_i_2, wb_dat_i_3, 
        wb_dat_i_4, wb_dat_i_5, wb_dat_i_6, wb_dat_i_7, wb_dat_i_8, wb_dat_i_9, 
        wb_dat_i_10, wb_dat_i_11, wb_dat_i_12, wb_dat_i_13, wb_dat_i_14, 
        wb_dat_i_15, wb_dat_i_16, wb_dat_i_17, wb_dat_i_18, wb_dat_i_19, 
        wb_dat_i_20, wb_dat_i_21, wb_dat_i_22, wb_dat_i_23, wb_dat_i_24, 
        wb_dat_i_25, wb_dat_i_26, wb_dat_i_27, wb_dat_i_28, wb_dat_i_29, 
        wb_dat_i_30, wb_dat_i_31, wb_adr_i_2, wb_adr_i_3, wb_adr_i_4, 
        wb_adr_i_5, wb_adr_i_6, wb_adr_i_7, wb_adr_i_8, wb_adr_i_9, 
        wb_adr_i_10, wb_adr_i_11, wb_sel_i_0, wb_sel_i_1, wb_sel_i_2, 
        wb_sel_i_3, m_wb_dat_i_0, m_wb_dat_i_1, m_wb_dat_i_2, m_wb_dat_i_3, 
        m_wb_dat_i_4, m_wb_dat_i_5, m_wb_dat_i_6, m_wb_dat_i_7, m_wb_dat_i_8, 
        m_wb_dat_i_9, m_wb_dat_i_10, m_wb_dat_i_11, m_wb_dat_i_12, 
        m_wb_dat_i_13, m_wb_dat_i_14, m_wb_dat_i_15, m_wb_dat_i_16, 
        m_wb_dat_i_17, m_wb_dat_i_18, m_wb_dat_i_19, m_wb_dat_i_20, 
        m_wb_dat_i_21, m_wb_dat_i_22, m_wb_dat_i_23, m_wb_dat_i_24, 
        m_wb_dat_i_25, m_wb_dat_i_26, m_wb_dat_i_27, m_wb_dat_i_28, 
        m_wb_dat_i_29, m_wb_dat_i_30, m_wb_dat_i_31, mrxd_pad_i_0, 
        mrxd_pad_i_1, mrxd_pad_i_2, mrxd_pad_i_3, wb_clk_i, wb_rst_i, wb_we_i, 
        wb_cyc_i, wb_stb_i, m_wb_ack_i, m_wb_err_i, mtx_clk_pad_i, 
        mrx_clk_pad_i, mrxdv_pad_i, mrxerr_pad_i, mcoll_pad_i, mcrs_pad_i, 
        md_pad_i, BD_WB_DAT_O_0, BD_WB_DAT_O_1, BD_WB_DAT_O_2, BD_WB_DAT_O_3, 
        BD_WB_DAT_O_4, BD_WB_DAT_O_5, BD_WB_DAT_O_6, BD_WB_DAT_O_7, 
        BD_WB_DAT_O_8, BD_WB_DAT_O_9, BD_WB_DAT_O_10, BD_WB_DAT_O_11, 
        BD_WB_DAT_O_12, BD_WB_DAT_O_13, BD_WB_DAT_O_14, BD_WB_DAT_O_15, 
        BD_WB_DAT_O_16, BD_WB_DAT_O_17, BD_WB_DAT_O_18, BD_WB_DAT_O_19, 
        BD_WB_DAT_O_20, BD_WB_DAT_O_21, BD_WB_DAT_O_22, BD_WB_DAT_O_23, 
        BD_WB_DAT_O_24, BD_WB_DAT_O_25, BD_WB_DAT_O_26, BD_WB_DAT_O_27, 
        BD_WB_DAT_O_28, BD_WB_DAT_O_29, BD_WB_DAT_O_30, BD_WB_DAT_O_31, 
        CarrierSense_Tx1, CarrierSense_Tx2, Collision_Tx1, RxAbortRst, 
        RxAbort_latch, RxAbort_sync1, RxAbort_wb, WillSendControlFrame_sync1, 
        WillSendControlFrame_sync2, WillSendControlFrame_sync3, RstTxPauseRq, 
        TxPauseRq_sync1, TxPauseRq_sync2, TxPauseRq_sync3, TPauseRq, RxEnSync, 
        Collision_Tx2, WillTransmit_q, WillTransmit_q2, p_miim1_LatchByte_0, 
        p_miim1_LatchByte0_d, p_miim1_LatchByte_1, p_miim1_LatchByte1_d, 
        p_miim1_WriteOp, p_miim1_BitCounter_6, p_miim1_BitCounter_4, 
        p_miim1_BitCounter_3, p_miim1_BitCounter_2, p_miim1_BitCounter_5, 
        p_miim1_BitCounter_1, NValid_stat, UpdateMIIRX_DATAReg, 
        p_miim1_WCtrlDataStart_q, p_miim1_RStatStart_q2, p_miim1_RStatStart_q1, 
        RStatStart, p_miim1_WCtrlDataStart_q2, p_miim1_WCtrlDataStart_q1, 
        WCtrlDataStart, p_miim1_EndBusy, p_miim1_InProgress_q3, 
        p_miim1_InProgress_q2, p_miim1_InProgress_q1, p_miim1_InProgress, 
        p_miim1_BitCounter_0, p_miim1_WCtrlData_q3, p_miim1_RStat_q3, 
        p_miim1_SyncStatMdcEn, p_miim1_ScanStat_q2, p_ethreg1_INT_SOURCEOut_6, 
        p_ethreg1_INT_SOURCEOut_5, p_ethreg1_INT_SOURCEOut_4, 
        p_ethreg1_INT_SOURCEOut_3, p_ethreg1_INT_SOURCEOut_2, 
        p_ethreg1_INT_SOURCEOut_1, p_ethreg1_INT_SOURCEOut_0, 
        p_ethreg1_SetRxCIrq, p_ethreg1_ResetRxCIrq_sync2, 
        p_ethreg1_SetRxCIrq_sync3, p_ethreg1_ResetRxCIrq_sync3, 
        p_ethreg1_SetTxCIrq, p_ethreg1_SetTxCIrq_sync3, 
        p_ethreg1_ResetTxCIrq_sync2, p_maccontrol1_MuxedDone, 
        p_maccontrol1_MuxedAbort, p_maccontrol1_TxDoneInLatched, 
        p_maccontrol1_TxAbortInLatched, p_maccontrol1_TxUsedDataOutDetected, 
        RetryCnt_2, RetryCnt_1, p_txethmac1_PacketFinished, TxRetry, 
        p_txethmac1_StatusLatch, p_txethmac1_ColWindow, 
        p_txethmac1_StopExcessiveDeferOccured, TxUsedDataIn, RetryCnt_3, 
        RetryCnt_0, p_txethmac1_PacketFinished_q, p_rxethmac1_Broadcast, 
        p_rxethmac1_Multicast, RxEndFrm, p_rxethmac1_RxEndFrm_d, RxStartFrm, 
        RxValid, RxData_7, RxData_6, RxData_5, RxData_4, RxData_3, RxData_2, 
        RxData_1, RxData_0, p_rxethmac1_DelayData, p_rxethmac1_LatchedByte_0, 
        p_rxethmac1_LatchedByte_1, p_rxethmac1_LatchedByte_2, 
        p_rxethmac1_LatchedByte_3, p_rxethmac1_CrcHash_0, 
        p_rxethmac1_CrcHash_1, p_rxethmac1_CrcHash_2, p_rxethmac1_CrcHash_3, 
        p_rxethmac1_CrcHash_4, p_rxethmac1_CrcHash_5, p_rxethmac1_CrcHashGood, 
        p_wishbone_Busy_IRQ_syncb1, p_wishbone_Busy_IRQ_sync3, 
        p_wishbone_Busy_IRQ_syncb2, RxE_IRQ, RxB_IRQ, TxE_IRQ, TxB_IRQ, 
        p_wishbone_RxStatusWriteLatched_syncb1, 
        p_wishbone_RxStatusWriteLatched_syncb2, p_wishbone_RxPointerMSB_30, 
        p_wishbone_RxPointerMSB_29, p_wishbone_RxPointerMSB_28, 
        p_wishbone_RxPointerMSB_27, p_wishbone_RxPointerMSB_26, 
        p_wishbone_RxPointerMSB_25, p_wishbone_RxPointerMSB_24, 
        p_wishbone_RxPointerMSB_23, p_wishbone_RxPointerMSB_22, 
        p_wishbone_RxPointerMSB_21, p_wishbone_RxPointerMSB_20, 
        p_wishbone_RxPointerMSB_19, p_wishbone_RxPointerMSB_18, 
        p_wishbone_RxPointerMSB_17, p_wishbone_RxPointerMSB_16, 
        p_wishbone_RxPointerMSB_15, p_wishbone_RxPointerMSB_14, 
        p_wishbone_RxPointerMSB_13, p_wishbone_RxPointerMSB_12, 
        p_wishbone_RxPointerMSB_11, p_wishbone_RxPointerMSB_10, 
        p_wishbone_RxPointerMSB_9, p_wishbone_RxPointerMSB_8, 
        p_wishbone_RxPointerMSB_7, p_wishbone_RxPointerMSB_6, 
        p_wishbone_RxPointerMSB_5, p_wishbone_RxPointerMSB_4, 
        p_wishbone_RxPointerMSB_3, p_wishbone_RxPointerMSB_2, 
        p_wishbone_RxPointerMSB_31, p_wishbone_TxPointerMSB_30, 
        p_wishbone_TxPointerMSB_29, p_wishbone_TxPointerMSB_28, 
        p_wishbone_TxPointerMSB_27, p_wishbone_TxPointerMSB_26, 
        p_wishbone_TxPointerMSB_25, p_wishbone_TxPointerMSB_24, 
        p_wishbone_TxPointerMSB_23, p_wishbone_TxPointerMSB_22, 
        p_wishbone_TxPointerMSB_21, p_wishbone_TxPointerMSB_20, 
        p_wishbone_TxPointerMSB_19, p_wishbone_TxPointerMSB_18, 
        p_wishbone_TxPointerMSB_17, p_wishbone_TxPointerMSB_16, 
        p_wishbone_TxPointerMSB_15, p_wishbone_TxPointerMSB_14, 
        p_wishbone_TxPointerMSB_13, p_wishbone_TxPointerMSB_12, 
        p_wishbone_TxPointerMSB_11, p_wishbone_TxPointerMSB_10, 
        p_wishbone_TxPointerMSB_9, p_wishbone_TxPointerMSB_8, 
        p_wishbone_TxPointerMSB_7, p_wishbone_TxPointerMSB_6, 
        p_wishbone_TxPointerMSB_5, p_wishbone_TxPointerMSB_4, 
        p_wishbone_TxPointerMSB_3, p_wishbone_TxPointerMSB_2, 
        p_wishbone_TxPointerMSB_31, p_wishbone_BlockingIncrementTxPointer, 
        p_wishbone_IncrTxPointer, p_wishbone_rx_burst_cnt_1, 
        p_wishbone_rx_burst_cnt_0, p_wishbone_TxAbortPacketBlocked, TxData_7, 
        p_wishbone_TxDataLatched_31, TxData_6, p_wishbone_TxDataLatched_30, 
        TxData_5, p_wishbone_TxDataLatched_29, TxData_4, 
        p_wishbone_TxDataLatched_28, TxData_3, p_wishbone_TxDataLatched_27, 
        TxData_2, p_wishbone_TxDataLatched_26, TxData_1, 
        p_wishbone_TxDataLatched_25, TxData_0, p_wishbone_TxDataLatched_24, 
        p_wishbone_TxDataLatched_23, p_wishbone_TxDataLatched_22, 
        p_wishbone_TxDataLatched_21, p_wishbone_TxDataLatched_20, 
        p_wishbone_TxDataLatched_19, p_wishbone_TxDataLatched_18, 
        p_wishbone_TxDataLatched_17, p_wishbone_TxDataLatched_16, 
        p_wishbone_TxDataLatched_15, p_wishbone_TxDataLatched_14, 
        p_wishbone_TxDataLatched_13, p_wishbone_TxDataLatched_12, 
        p_wishbone_TxDataLatched_11, p_wishbone_TxDataLatched_10, 
        p_wishbone_TxDataLatched_9, p_wishbone_TxDataLatched_8, 
        p_wishbone_TxDataLatched_7, p_wishbone_TxDataLatched_6, 
        p_wishbone_TxDataLatched_5, p_wishbone_TxDataLatched_4, 
        p_wishbone_TxDataLatched_3, p_wishbone_TxDataLatched_2, 
        p_wishbone_TxDataLatched_1, p_wishbone_TxDataLatched_0, 
        p_wishbone_StartOccured, p_wishbone_TxByteCnt_1, 
        p_wishbone_TxByteCnt_0, TxStartFrm, p_wishbone_TxStartFrm_syncb2, 
        p_wishbone_TxEndFrm_wb, p_wishbone_ram_di_8, TxUnderRun, 
        p_wishbone_TxUnderRun_sync1, p_wishbone_TxUnderRun_wb, 
        p_wishbone_TxAbortPacket, p_wishbone_BlockingTxStatusWrite_sync3, 
        p_wishbone_ram_addr_1, p_wishbone_ram_addr_7, p_wishbone_TxBDAddress_7, 
        p_wishbone_ram_addr_6, p_wishbone_TxBDAddress_6, p_wishbone_ram_addr_5, 
        p_wishbone_TxBDAddress_5, p_wishbone_ram_addr_4, 
        p_wishbone_TxBDAddress_4, p_wishbone_ram_addr_3, 
        p_wishbone_TxBDAddress_3, p_wishbone_ram_addr_2, 
        p_wishbone_TxBDAddress_2, p_wishbone_TxBDAddress_1, 
        p_wishbone_TxRetryPacket_NotCleared, p_wishbone_ram_addr_0, 
        p_wishbone_TxPointerLSB_1, p_wishbone_TxPointerLSB_0, 
        p_wishbone_ram_di_14, p_wishbone_ram_di_15, p_wishbone_ram_di_10, 
        p_wishbone_ram_di_9, BDAck, p_wishbone_BDRead, p_wishbone_ram_di_31, 
        p_wishbone_ram_di_30, p_wishbone_ram_di_29, p_wishbone_ram_di_28, 
        p_wishbone_ram_di_27, p_wishbone_ram_di_26, p_wishbone_ram_di_25, 
        p_wishbone_ram_di_24, p_wishbone_ram_di_23, p_wishbone_ram_di_22, 
        p_wishbone_ram_di_21, p_wishbone_ram_di_20, p_wishbone_ram_di_19, 
        p_wishbone_ram_di_18, p_wishbone_ram_di_17, p_wishbone_ram_di_16, 
        p_wishbone_ram_di_13, p_wishbone_ram_di_12, p_wishbone_ram_di_11, 
        p_wishbone_ram_di_7, p_wishbone_ram_di_5, p_wishbone_ram_di_4, 
        p_wishbone_ram_di_3, p_wishbone_ram_di_2, p_wishbone_ram_di_1, 
        p_wishbone_ram_di_0, p_wishbone_BDWrite_0, p_wishbone_BDWrite_1, 
        p_wishbone_BDWrite_2, p_wishbone_BDWrite_3, p_wishbone_RxBDDataIn_14, 
        p_wishbone_RxBDAddress_7, p_wishbone_RxBDAddress_6, 
        p_wishbone_RxBDAddress_5, p_wishbone_RxBDAddress_4, 
        p_wishbone_RxBDAddress_3, p_wishbone_RxBDAddress_2, 
        p_wishbone_RxBDAddress_1, p_wishbone_RxBDDataIn_13, 
        p_wishbone_ShiftEndedSync3, p_wishbone_RxDataLatched2_8, 
        p_wishbone_RxDataLatched1_8, p_wishbone_RxDataLatched2_9, 
        p_wishbone_RxDataLatched1_9, p_wishbone_RxDataLatched2_10, 
        p_wishbone_RxDataLatched1_10, p_wishbone_RxDataLatched2_11, 
        p_wishbone_RxDataLatched1_11, p_wishbone_RxDataLatched2_12, 
        p_wishbone_RxDataLatched1_12, p_wishbone_RxDataLatched2_13, 
        p_wishbone_RxDataLatched1_13, p_wishbone_RxDataLatched2_14, 
        p_wishbone_RxDataLatched1_14, p_wishbone_RxDataLatched2_15, 
        p_wishbone_RxDataLatched1_15, p_wishbone_RxDataLatched2_24, 
        p_wishbone_RxDataLatched1_24, p_wishbone_RxDataLatched2_25, 
        p_wishbone_RxDataLatched1_25, p_wishbone_RxDataLatched2_26, 
        p_wishbone_RxDataLatched1_26, p_wishbone_RxDataLatched2_27, 
        p_wishbone_RxDataLatched1_27, p_wishbone_RxDataLatched2_28, 
        p_wishbone_RxDataLatched1_28, p_wishbone_RxDataLatched2_29, 
        p_wishbone_RxDataLatched1_29, p_wishbone_RxDataLatched2_30, 
        p_wishbone_RxDataLatched1_30, p_wishbone_RxDataLatched2_31, 
        p_wishbone_RxDataLatched1_31, p_wishbone_RxDataLatched2_17, 
        p_wishbone_RxDataLatched2_18, p_wishbone_RxDataLatched2_19, 
        p_wishbone_RxDataLatched2_20, p_wishbone_RxDataLatched2_21, 
        p_wishbone_RxDataLatched2_22, p_wishbone_RxDataLatched2_23, 
        p_wishbone_RxDataLatched2_0, p_wishbone_RxDataLatched2_1, 
        p_wishbone_RxDataLatched2_2, p_wishbone_RxDataLatched2_3, 
        p_wishbone_RxDataLatched2_4, p_wishbone_RxDataLatched2_5, 
        p_wishbone_RxDataLatched2_6, p_wishbone_RxDataLatched2_7, 
        p_wishbone_WriteRxDataToFifoSync3, p_wishbone_RxByteCnt_1, 
        p_wishbone_RxByteCnt_0, p_wishbone_ShiftWillEnd, 
        p_wishbone_ShiftEndedSync_c2, p_wishbone_RxValidBytes_1, 
        p_wishbone_RxValidBytes_0, p_wishbone_LastByteIn, p_wishbone_RxBDRead, 
        p_wishbone_RxReady, p_wishbone_ShiftEnded, 
        p_wishbone_RxDataLatched2_16, p_wishbone_RxDataLatched1_16, 
        p_wishbone_RxDataLatched1_17, p_wishbone_RxDataLatched1_18, 
        p_wishbone_RxDataLatched1_19, p_wishbone_RxDataLatched1_20, 
        p_wishbone_RxDataLatched1_21, p_wishbone_RxDataLatched1_22, 
        p_wishbone_RxDataLatched1_23, p_wishbone_RxPointerLSB_rst_0, 
        p_wishbone_RxPointerLSB_rst_1, p_wishbone_RxPointerRead, 
        p_wishbone_RxBDReady, p_wishbone_RxEn_q, p_wishbone_RxEn_needed, 
        p_wishbone_WbEn_q, p_wishbone_LatchedTxLength_15, 
        p_wishbone_LatchedTxLength_14, p_wishbone_LatchedTxLength_13, 
        p_wishbone_LatchedTxLength_12, p_wishbone_LatchedTxLength_11, 
        p_wishbone_LatchedTxLength_10, p_wishbone_LatchedTxLength_9, 
        p_wishbone_LatchedTxLength_8, p_wishbone_LatchedTxLength_7, 
        p_wishbone_LatchedTxLength_6, p_wishbone_LatchedTxLength_5, 
        p_wishbone_LatchedTxLength_4, p_wishbone_LatchedTxLength_3, 
        p_wishbone_LatchedTxLength_2, p_wishbone_LatchedTxLength_1, 
        p_wishbone_LatchedTxLength_0, p_wishbone_BlockingTxBDRead, 
        p_wishbone_TxBDReady, p_wishbone_ReadTxDataFromMemory, 
        p_wishbone_TxLength_14, p_wishbone_TxLength_13, p_wishbone_TxLength_12, 
        p_wishbone_TxLength_11, p_wishbone_TxLength_10, p_wishbone_TxLength_9, 
        p_wishbone_TxLength_8, p_wishbone_TxLength_7, p_wishbone_TxLength_6, 
        p_wishbone_TxLength_5, p_wishbone_TxLength_4, p_wishbone_TxLength_3, 
        p_wishbone_TxLength_2, p_wishbone_TxValidBytesLatched_1, 
        p_wishbone_TxLength_1, p_wishbone_TxLength_0, PerPacketCrcEn, 
        PerPacketPad, p_wishbone_TxStatus_13, p_wishbone_TxStatus_14, 
        p_wishbone_TxDonePacket_NotCleared, p_wishbone_TxEn_q, 
        p_wishbone_TxEn_needed, p_wishbone_U3_U3_Z_0, 
        p_wishbone_TxPointerLSB_rst_1, p_wishbone_TxPointerRead, 
        p_wishbone_TxBDRead, p_wishbone_TxAbortPacket_NotCleared, 
        p_wishbone_TxRetryPacketBlocked, p_wishbone_TxRetryPacket, 
        p_wishbone_TxDonePacketBlocked, p_wishbone_TxDonePacket, 
        p_wishbone_tx_burst_en, p_wishbone_tx_burst_cnt_2, 
        p_wishbone_tx_burst_cnt_1, p_wishbone_tx_burst_cnt_0, 
        p_wishbone_cyc_cleared, p_wishbone_MasterWbTX, p_wishbone_MasterWbRX, 
        p_wishbone_rx_burst_en, p_wishbone_rx_burst_cnt_2, 
        p_wishbone_BlockReadTxDataFromMemory, 
        p_wishbone_ReadTxDataFromFifo_sync3, 
        p_wishbone_ReadTxDataFromFifo_syncb3, p_wishbone_LastWord, TxEndFrm, 
        p_wishbone_TxValidBytesLatched_0, p_wishbone_LatchValidBytes_q, 
        p_wishbone_TxLength_15, p_wishbone_ram_di_6, p_wishbone_RxBDDataIn_6, 
        p_wishbone_RxStatusIn_6, p_wishbone_RxBDDataIn_0, 
        p_wishbone_RxBDDataIn_1, p_wishbone_RxBDDataIn_2, 
        p_wishbone_RxBDDataIn_3, p_wishbone_RxBDDataIn_4, 
        p_wishbone_RxBDDataIn_5, p_wishbone_RxBDDataIn_7, 
        p_wishbone_RxBDDataIn_8, p_wishbone_RxBDDataIn_16, 
        p_wishbone_RxBDDataIn_17, p_wishbone_RxBDDataIn_18, 
        p_wishbone_RxBDDataIn_19, p_wishbone_RxBDDataIn_20, 
        p_wishbone_RxBDDataIn_21, p_wishbone_RxBDDataIn_22, 
        p_wishbone_RxBDDataIn_23, p_wishbone_RxBDDataIn_24, 
        p_wishbone_RxBDDataIn_25, p_wishbone_RxBDDataIn_26, 
        p_wishbone_RxBDDataIn_27, p_wishbone_RxBDDataIn_28, 
        p_wishbone_RxBDDataIn_29, p_wishbone_RxBDDataIn_30, 
        p_wishbone_RxBDDataIn_31, p_wishbone_RxAbortSyncb2, 
        p_wishbone_RxAbortSync4, p_wishbone_RxEnableWindow, 
        p_wishbone_SyncRxStartFrm_q2, p_wishbone_SyncRxStartFrm, 
        p_wishbone_TxAbort_wb_q, p_wishbone_TxDone_wb_q, 
        p_wishbone_TxRetry_wb_q, p_wishbone_TxAbort_q, p_wishbone_TxUsedData_q, 
        p_wishbone_Flop, p_wishbone_TxRetry_q, p_wishbone_r_RxEn_q, 
        p_wishbone_r_TxEn_q, CarrierSenseLost, DeferLatched, LateCollLatched, 
        RetryLimit, RetryCntLatched_0, RetryCntLatched_1, RetryCntLatched_2, 
        RetryCntLatched_3, ReceivedPacketTooBig, DribbleNibble, ShortFrame, 
        RxLateCollision, p_macstatus1_RxColWindow, InvalidSymbol, ReceiveEnd, 
        LatchedMRxErr, LatchedCrcError, p_miim1_clkgen_Counter_6, 
        p_miim1_clkgen_Counter_5, p_miim1_clkgen_Counter_4, 
        p_miim1_clkgen_Counter_3, p_miim1_clkgen_Counter_2, 
        p_miim1_clkgen_Counter_1, p_miim1_clkgen_Counter_0, LinkFail, Prsd_0, 
        Prsd_1, Prsd_2, Prsd_3, Prsd_4, Prsd_5, Prsd_6, Prsd_7, Prsd_8, Prsd_9, 
        Prsd_10, Prsd_11, Prsd_12, Prsd_13, Prsd_14, Prsd_15, 
        p_miim1_ShiftedBit, p_miim1_shftrg_ShiftReg_6, 
        p_miim1_shftrg_ShiftReg_5, p_miim1_shftrg_ShiftReg_4, 
        p_miim1_shftrg_ShiftReg_3, p_miim1_shftrg_ShiftReg_2, 
        p_miim1_shftrg_ShiftReg_1, p_miim1_shftrg_ShiftReg_0, 
        p_miim1_outctrl_Mdo_d, p_miim1_outctrl_Mdo_2d, p_miim1_outctrl_MdoEn_d, 
        p_miim1_outctrl_MdoEn_2d, p_ethreg1_MODEROut_0, p_ethreg1_MODEROut_1, 
        p_ethreg1_r_NoPre, r_Bro, p_ethreg1_r_Iam, r_Pro, r_IFG, r_LoopBck, 
        r_NoBckof, r_ExDfrEn, r_FullD, p_ethreg1_MODEROut_11, r_DlyCrcEn, 
        r_CrcEn, r_HugEn, r_Pad, r_RecSmall, p_ethreg1_INT_MASKOut_0, 
        p_ethreg1_INT_MASKOut_1, p_ethreg1_INT_MASKOut_2, 
        p_ethreg1_INT_MASKOut_3, p_ethreg1_INT_MASKOut_4, 
        p_ethreg1_INT_MASKOut_5, p_ethreg1_INT_MASKOut_6, r_IPGT_0, r_IPGT_1, 
        r_IPGT_2, r_IPGT_3, r_IPGT_4, r_IPGT_5, r_IPGT_6, r_IPGR1_0, r_IPGR1_1, 
        r_IPGR1_2, r_IPGR1_3, r_IPGR1_4, r_IPGR1_5, r_IPGR1_6, r_MaxFL_8, 
        r_MaxFL_9, r_MaxFL_10, r_MaxFL_11, r_MaxFL_12, r_MaxFL_13, r_MaxFL_14, 
        r_MaxFL_15, p_txethmac1_txcounters1_N41, p_txethmac1_txcounters1_N42, 
        r_MinFL_2, r_MinFL_3, r_MinFL_4, r_MinFL_5, r_MinFL_6, r_MinFL_7, 
        r_CollValid_0, r_CollValid_1, r_CollValid_2, r_CollValid_3, 
        r_CollValid_4, r_CollValid_5, r_MaxRet_0, r_MaxRet_1, r_MaxRet_2, 
        r_MaxRet_3, r_PassAll, r_RxFlow, r_TxFlow, r_ClkDiv_0, r_ClkDiv_1, 
        r_ClkDiv_2, r_ClkDiv_3, r_ClkDiv_4, r_ClkDiv_5, r_ClkDiv_6, r_ClkDiv_7, 
        r_FIAD_0, r_FIAD_1, r_FIAD_2, r_FIAD_3, r_FIAD_4, 
        p_ethreg1_MIIRX_DATAOut_0, p_ethreg1_MIIRX_DATAOut_1, 
        p_ethreg1_MIIRX_DATAOut_2, p_ethreg1_MIIRX_DATAOut_3, 
        p_ethreg1_MIIRX_DATAOut_4, p_ethreg1_MIIRX_DATAOut_5, 
        p_ethreg1_MIIRX_DATAOut_6, p_ethreg1_MIIRX_DATAOut_7, 
        p_ethreg1_MIIRX_DATAOut_8, p_ethreg1_MIIRX_DATAOut_9, 
        p_ethreg1_MIIRX_DATAOut_10, p_ethreg1_MIIRX_DATAOut_11, 
        p_ethreg1_MIIRX_DATAOut_12, p_ethreg1_MIIRX_DATAOut_13, 
        p_ethreg1_MIIRX_DATAOut_14, p_ethreg1_MIIRX_DATAOut_15, 
        ReceivedPauseFrm, p_maccontrol1_receivecontrol1_SlotTimer_4, 
        p_maccontrol1_receivecontrol1_SlotTimer_3, 
        p_maccontrol1_receivecontrol1_SlotTimer_2, 
        p_maccontrol1_receivecontrol1_SlotTimer_1, 
        p_maccontrol1_receivecontrol1_SlotTimer_5, p_maccontrol1_Pause, 
        p_maccontrol1_receivecontrol1_PauseTimerEq0_sync2, 
        p_maccontrol1_receivecontrol1_Divider2, 
        p_maccontrol1_receivecontrol1_PauseTimer_15, 
        p_maccontrol1_receivecontrol1_PauseTimer_14, 
        p_maccontrol1_receivecontrol1_PauseTimer_13, 
        p_maccontrol1_receivecontrol1_PauseTimer_12, 
        p_maccontrol1_receivecontrol1_PauseTimer_11, 
        p_maccontrol1_receivecontrol1_PauseTimer_10, 
        p_maccontrol1_receivecontrol1_PauseTimer_9, 
        p_maccontrol1_receivecontrol1_PauseTimer_8, 
        p_maccontrol1_receivecontrol1_PauseTimer_7, 
        p_maccontrol1_receivecontrol1_PauseTimer_6, 
        p_maccontrol1_receivecontrol1_PauseTimer_5, 
        p_maccontrol1_receivecontrol1_PauseTimer_4, 
        p_maccontrol1_receivecontrol1_PauseTimer_3, 
        p_maccontrol1_receivecontrol1_PauseTimer_2, 
        p_maccontrol1_receivecontrol1_PauseTimer_1, 
        p_maccontrol1_receivecontrol1_PauseTimer_0, 
        p_maccontrol1_receivecontrol1_SlotTimer_0, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_0, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_1, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_2, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_3, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_4, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_5, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_6, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_7, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_8, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_9, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_10, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_11, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_12, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_13, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_14, 
        p_maccontrol1_receivecontrol1_LatchedTimerValue_15, 
        p_maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr, 
        ControlFrmAddressOK, p_maccontrol1_receivecontrol1_OpCodeOK, 
        p_maccontrol1_receivecontrol1_TypeLengthOK, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_0, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_1, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_2, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_3, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_4, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_5, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_6, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_7, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_8, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_9, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_10, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_11, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_12, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_13, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_14, 
        p_maccontrol1_receivecontrol1_AssembledTimerValue_15, 
        p_maccontrol1_receivecontrol1_ByteCnt_3, 
        p_maccontrol1_receivecontrol1_ByteCnt_2, 
        p_maccontrol1_receivecontrol1_ByteCnt_1, 
        p_maccontrol1_receivecontrol1_ByteCnt_4, 
        p_maccontrol1_receivecontrol1_DetectionWindow, 
        p_maccontrol1_receivecontrol1_ByteCnt_0, 
        p_maccontrol1_receivecontrol1_DlyCrcCnt_1, 
        p_maccontrol1_receivecontrol1_DlyCrcCnt_2, 
        p_maccontrol1_receivecontrol1_DlyCrcCnt_0, p_maccontrol1_ControlData_0, 
        p_maccontrol1_ControlData_1, p_maccontrol1_ControlData_2, 
        p_maccontrol1_ControlData_3, p_maccontrol1_ControlData_4, 
        p_maccontrol1_ControlData_5, p_maccontrol1_ControlData_6, 
        p_maccontrol1_ControlData_7, p_maccontrol1_transmitcontrol1_ByteCnt_4, 
        p_maccontrol1_transmitcontrol1_ByteCnt_3, 
        p_maccontrol1_transmitcontrol1_ByteCnt_2, 
        p_maccontrol1_transmitcontrol1_ByteCnt_1, 
        p_maccontrol1_transmitcontrol1_ByteCnt_5, 
        p_maccontrol1_transmitcontrol1_DlyCrcCnt_2, 
        p_maccontrol1_transmitcontrol1_DlyCrcCnt_1, 
        p_maccontrol1_transmitcontrol1_DlyCrcCnt_0, p_maccontrol1_BlockTxDone, 
        p_maccontrol1_SendingCtrlFrm, 
        p_maccontrol1_transmitcontrol1_TxCtrlStartFrm_q, p_maccontrol1_CtrlMux, 
        TxCtrlEndFrm, p_maccontrol1_transmitcontrol1_ControlEnd_q, 
        p_maccontrol1_transmitcontrol1_ByteCnt_0, 
        p_maccontrol1_transmitcontrol1_TxUsedDataIn_q, p_txethmac1_DlyCrcCnt_1, 
        p_txethmac1_DlyCrcCnt_2, p_txethmac1_DlyCrcCnt_0, 
        p_txethmac1_txcounters1_ByteCnt_14, p_txethmac1_txcounters1_ByteCnt_13, 
        p_txethmac1_txcounters1_ByteCnt_12, p_txethmac1_txcounters1_ByteCnt_11, 
        p_txethmac1_txcounters1_ByteCnt_10, p_txethmac1_ByteCnt_9, 
        p_txethmac1_ByteCnt_8, p_txethmac1_ByteCnt_7, p_txethmac1_ByteCnt_6, 
        p_txethmac1_ByteCnt_5, p_txethmac1_ByteCnt_4, p_txethmac1_ByteCnt_3, 
        p_txethmac1_ByteCnt_2, p_txethmac1_ByteCnt_1, 
        p_txethmac1_txcounters1_ByteCnt_15, p_txethmac1_ByteCnt_0, 
        p_txethmac1_NibCnt_15, p_txethmac1_NibCnt_14, p_txethmac1_NibCnt_13, 
        p_txethmac1_NibCnt_12, p_txethmac1_NibCnt_11, p_txethmac1_NibCnt_10, 
        p_txethmac1_NibCnt_9, p_txethmac1_NibCnt_8, p_txethmac1_NibCnt_7, 
        p_txethmac1_NibCnt_6, p_txethmac1_NibCnt_5, p_txethmac1_NibCnt_4, 
        p_txethmac1_NibCnt_2, p_txethmac1_NibCnt_1, p_txethmac1_NibCnt_3, 
        p_txethmac1_NibCnt_0, p_txethmac1_StateBackOff, p_txethmac1_StateJam_q, 
        p_txethmac1_StatePAD, StateData_1, StateData_0, StatePreamble, 
        p_txethmac1_StateFCS, p_txethmac1_StateIdle, p_txethmac1_StateDefer, 
        p_txethmac1_StateIPG, p_txethmac1_txstatem1_Rule1, 
        p_txethmac1_txcrc_Crc_22, p_txethmac1_txcrc_Crc_18, 
        p_txethmac1_txcrc_Crc_14, p_txethmac1_txcrc_Crc_10, 
        p_txethmac1_txcrc_Crc_6, p_txethmac1_txcrc_Crc_2, 
        p_txethmac1_txcrc_Crc_5, p_txethmac1_txcrc_Crc_23, 
        p_txethmac1_txcrc_Crc_19, p_txethmac1_txcrc_Crc_15, 
        p_txethmac1_txcrc_Crc_11, p_txethmac1_txcrc_Crc_7, 
        p_txethmac1_txcrc_Crc_3, p_txethmac1_Crc_31, p_txethmac1_txcrc_Crc_27, 
        p_txethmac1_txcrc_Crc_1, p_txethmac1_Crc_29, p_txethmac1_txcrc_Crc_25, 
        p_txethmac1_txcrc_Crc_21, p_txethmac1_txcrc_Crc_17, 
        p_txethmac1_txcrc_Crc_13, p_txethmac1_txcrc_Crc_9, p_txethmac1_Crc_30, 
        p_txethmac1_txcrc_Crc_26, p_txethmac1_Crc_28, p_txethmac1_txcrc_Crc_24, 
        p_txethmac1_txcrc_Crc_20, p_txethmac1_txcrc_Crc_16, 
        p_txethmac1_txcrc_Crc_12, p_txethmac1_txcrc_Crc_8, 
        p_txethmac1_txcrc_Crc_4, p_txethmac1_txcrc_Crc_0, 
        p_txethmac1_random1_RandomLatched_0, 
        p_txethmac1_random1_RandomLatched_1, 
        p_txethmac1_random1_RandomLatched_2, 
        p_txethmac1_random1_RandomLatched_3, 
        p_txethmac1_random1_RandomLatched_4, 
        p_txethmac1_random1_RandomLatched_5, 
        p_txethmac1_random1_RandomLatched_6, 
        p_txethmac1_random1_RandomLatched_7, 
        p_txethmac1_random1_RandomLatched_8, 
        p_txethmac1_random1_RandomLatched_9, p_txethmac1_random1_x_9, 
        RxStateSFD, RxStateData_1, RxStatePreamble, RxStateIdle, 
        p_rxethmac1_StateDrop, p_rxethmac1_rxcounters1_ByteCnt_14, 
        p_rxethmac1_rxcounters1_ByteCnt_13, p_rxethmac1_rxcounters1_ByteCnt_12, 
        p_rxethmac1_rxcounters1_ByteCnt_11, p_rxethmac1_rxcounters1_ByteCnt_10, 
        p_rxethmac1_rxcounters1_ByteCnt_9, p_rxethmac1_rxcounters1_ByteCnt_8, 
        p_rxethmac1_rxcounters1_ByteCnt_7, p_rxethmac1_rxcounters1_ByteCnt_6, 
        p_rxethmac1_rxcounters1_ByteCnt_5, p_rxethmac1_rxcounters1_ByteCnt_4, 
        p_rxethmac1_rxcounters1_ByteCnt_3, p_rxethmac1_rxcounters1_ByteCnt_2, 
        RxByteCnt_1, p_rxethmac1_rxcounters1_ByteCnt_15, RxByteCnt_0, 
        p_rxethmac1_DlyCrcCnt_2, p_rxethmac1_DlyCrcCnt_1, 
        p_rxethmac1_DlyCrcCnt_3, p_rxethmac1_DlyCrcCnt_0, 
        p_rxethmac1_rxcounters1_IFGCounter_3, 
        p_rxethmac1_rxcounters1_IFGCounter_2, 
        p_rxethmac1_rxcounters1_IFGCounter_1, 
        p_rxethmac1_rxcounters1_IFGCounter_4, 
        p_rxethmac1_rxcounters1_IFGCounter_0, AddressMiss, 
        p_rxethmac1_rxaddrcheck1_MulticastOK, RxAbort, 
        p_rxethmac1_rxaddrcheck1_UnicastOK, p_wishbone_bd_ram_mem2_0_16, 
        p_wishbone_bd_ram_mem2_0_17, p_wishbone_bd_ram_mem2_0_18, 
        p_wishbone_bd_ram_mem2_0_19, p_wishbone_bd_ram_mem2_0_20, 
        p_wishbone_bd_ram_mem2_0_21, p_wishbone_bd_ram_mem2_0_22, 
        p_wishbone_bd_ram_mem2_0_23, p_wishbone_bd_ram_mem2_1_16, 
        p_wishbone_bd_ram_mem2_1_17, p_wishbone_bd_ram_mem2_1_18, 
        p_wishbone_bd_ram_mem2_1_19, p_wishbone_bd_ram_mem2_1_20, 
        p_wishbone_bd_ram_mem2_1_21, p_wishbone_bd_ram_mem2_1_22, 
        p_wishbone_bd_ram_mem2_1_23, p_wishbone_bd_ram_mem2_2_16, 
        p_wishbone_bd_ram_mem2_2_17, p_wishbone_bd_ram_mem2_2_18, 
        p_wishbone_bd_ram_mem2_2_19, p_wishbone_bd_ram_mem2_2_20, 
        p_wishbone_bd_ram_mem2_2_21, p_wishbone_bd_ram_mem2_2_22, 
        p_wishbone_bd_ram_mem2_2_23, p_wishbone_bd_ram_mem2_3_16, 
        p_wishbone_bd_ram_mem2_3_17, p_wishbone_bd_ram_mem2_3_18, 
        p_wishbone_bd_ram_mem2_3_19, p_wishbone_bd_ram_mem2_3_20, 
        p_wishbone_bd_ram_mem2_3_21, p_wishbone_bd_ram_mem2_3_22, 
        p_wishbone_bd_ram_mem2_3_23, p_wishbone_bd_ram_mem2_4_16, 
        p_wishbone_bd_ram_mem2_4_17, p_wishbone_bd_ram_mem2_4_18, 
        p_wishbone_bd_ram_mem2_4_19, p_wishbone_bd_ram_mem2_4_20, 
        p_wishbone_bd_ram_mem2_4_21, p_wishbone_bd_ram_mem2_4_22, 
        p_wishbone_bd_ram_mem2_4_23, p_wishbone_bd_ram_mem2_5_16, 
        p_wishbone_bd_ram_mem2_5_17, p_wishbone_bd_ram_mem2_5_18, 
        p_wishbone_bd_ram_mem2_5_19, p_wishbone_bd_ram_mem2_5_20, 
        p_wishbone_bd_ram_mem2_5_21, p_wishbone_bd_ram_mem2_5_22, 
        p_wishbone_bd_ram_mem2_5_23, p_wishbone_bd_ram_mem2_6_16, 
        p_wishbone_bd_ram_mem2_6_17, p_wishbone_bd_ram_mem2_6_18, 
        p_wishbone_bd_ram_mem2_6_19, p_wishbone_bd_ram_mem2_6_20, 
        p_wishbone_bd_ram_mem2_6_21, p_wishbone_bd_ram_mem2_6_22, 
        p_wishbone_bd_ram_mem2_6_23, p_wishbone_bd_ram_mem2_7_16, 
        p_wishbone_bd_ram_mem2_7_17, p_wishbone_bd_ram_mem2_7_18, 
        p_wishbone_bd_ram_mem2_7_19, p_wishbone_bd_ram_mem2_7_20, 
        p_wishbone_bd_ram_mem2_7_21, p_wishbone_bd_ram_mem2_7_22, 
        p_wishbone_bd_ram_mem2_7_23, p_wishbone_bd_ram_mem2_8_16, 
        p_wishbone_bd_ram_mem2_8_17, p_wishbone_bd_ram_mem2_8_18, 
        p_wishbone_bd_ram_mem2_8_19, p_wishbone_bd_ram_mem2_8_20, 
        p_wishbone_bd_ram_mem2_8_21, p_wishbone_bd_ram_mem2_8_22, 
        p_wishbone_bd_ram_mem2_8_23, p_wishbone_bd_ram_mem2_9_16, 
        p_wishbone_bd_ram_mem2_9_17, p_wishbone_bd_ram_mem2_9_18, 
        p_wishbone_bd_ram_mem2_9_19, p_wishbone_bd_ram_mem2_9_20, 
        p_wishbone_bd_ram_mem2_9_21, p_wishbone_bd_ram_mem2_9_22, 
        p_wishbone_bd_ram_mem2_9_23, p_wishbone_bd_ram_mem2_10_16, 
        p_wishbone_bd_ram_mem2_10_17, p_wishbone_bd_ram_mem2_10_18, 
        p_wishbone_bd_ram_mem2_10_19, p_wishbone_bd_ram_mem2_10_20, 
        p_wishbone_bd_ram_mem2_10_21, p_wishbone_bd_ram_mem2_10_22, 
        p_wishbone_bd_ram_mem2_10_23, p_wishbone_bd_ram_mem2_11_16, 
        p_wishbone_bd_ram_mem2_11_17, p_wishbone_bd_ram_mem2_11_18, 
        p_wishbone_bd_ram_mem2_11_19, p_wishbone_bd_ram_mem2_11_20, 
        p_wishbone_bd_ram_mem2_11_21, p_wishbone_bd_ram_mem2_11_22, 
        p_wishbone_bd_ram_mem2_11_23, p_wishbone_bd_ram_mem2_12_16, 
        p_wishbone_bd_ram_mem2_12_17, p_wishbone_bd_ram_mem2_12_18, 
        p_wishbone_bd_ram_mem2_12_19, p_wishbone_bd_ram_mem2_12_20, 
        p_wishbone_bd_ram_mem2_12_21, p_wishbone_bd_ram_mem2_12_22, 
        p_wishbone_bd_ram_mem2_12_23, p_wishbone_bd_ram_mem2_13_16, 
        p_wishbone_bd_ram_mem2_13_17, p_wishbone_bd_ram_mem2_13_18, 
        p_wishbone_bd_ram_mem2_13_19, p_wishbone_bd_ram_mem2_13_20, 
        p_wishbone_bd_ram_mem2_13_21, p_wishbone_bd_ram_mem2_13_22, 
        p_wishbone_bd_ram_mem2_13_23, p_wishbone_bd_ram_mem2_14_16, 
        p_wishbone_bd_ram_mem2_14_17, p_wishbone_bd_ram_mem2_14_18, 
        p_wishbone_bd_ram_mem2_14_19, p_wishbone_bd_ram_mem2_14_20, 
        p_wishbone_bd_ram_mem2_14_21, p_wishbone_bd_ram_mem2_14_22, 
        p_wishbone_bd_ram_mem2_14_23, p_wishbone_bd_ram_mem2_15_16, 
        p_wishbone_bd_ram_mem2_15_17, p_wishbone_bd_ram_mem2_15_18, 
        p_wishbone_bd_ram_mem2_15_19, p_wishbone_bd_ram_mem2_15_20, 
        p_wishbone_bd_ram_mem2_15_21, p_wishbone_bd_ram_mem2_15_22, 
        p_wishbone_bd_ram_mem2_15_23, p_wishbone_bd_ram_mem2_16_16, 
        p_wishbone_bd_ram_mem2_16_17, p_wishbone_bd_ram_mem2_16_18, 
        p_wishbone_bd_ram_mem2_16_19, p_wishbone_bd_ram_mem2_16_20, 
        p_wishbone_bd_ram_mem2_16_21, p_wishbone_bd_ram_mem2_16_22, 
        p_wishbone_bd_ram_mem2_16_23, p_wishbone_bd_ram_mem2_17_16, 
        p_wishbone_bd_ram_mem2_17_17, p_wishbone_bd_ram_mem2_17_18, 
        p_wishbone_bd_ram_mem2_17_19, p_wishbone_bd_ram_mem2_17_20, 
        p_wishbone_bd_ram_mem2_17_21, p_wishbone_bd_ram_mem2_17_22, 
        p_wishbone_bd_ram_mem2_17_23, p_wishbone_bd_ram_mem2_18_16, 
        p_wishbone_bd_ram_mem2_18_17, p_wishbone_bd_ram_mem2_18_18, 
        p_wishbone_bd_ram_mem2_18_19, p_wishbone_bd_ram_mem2_18_20, 
        p_wishbone_bd_ram_mem2_18_21, p_wishbone_bd_ram_mem2_18_22, 
        p_wishbone_bd_ram_mem2_18_23, p_wishbone_bd_ram_mem2_19_16, 
        p_wishbone_bd_ram_mem2_19_17, p_wishbone_bd_ram_mem2_19_18, 
        p_wishbone_bd_ram_mem2_19_19, p_wishbone_bd_ram_mem2_19_20, 
        p_wishbone_bd_ram_mem2_19_21, p_wishbone_bd_ram_mem2_19_22, 
        p_wishbone_bd_ram_mem2_19_23, p_wishbone_bd_ram_mem2_20_16, 
        p_wishbone_bd_ram_mem2_20_17, p_wishbone_bd_ram_mem2_20_18, 
        p_wishbone_bd_ram_mem2_20_19, p_wishbone_bd_ram_mem2_20_20, 
        p_wishbone_bd_ram_mem2_20_21, p_wishbone_bd_ram_mem2_20_22, 
        p_wishbone_bd_ram_mem2_20_23, p_wishbone_bd_ram_mem2_21_16, 
        p_wishbone_bd_ram_mem2_21_17, p_wishbone_bd_ram_mem2_21_18, 
        p_wishbone_bd_ram_mem2_21_19, p_wishbone_bd_ram_mem2_21_20, 
        p_wishbone_bd_ram_mem2_21_21, p_wishbone_bd_ram_mem2_21_22, 
        p_wishbone_bd_ram_mem2_21_23, p_wishbone_bd_ram_mem2_22_16, 
        p_wishbone_bd_ram_mem2_22_17, p_wishbone_bd_ram_mem2_22_18, 
        p_wishbone_bd_ram_mem2_22_19, p_wishbone_bd_ram_mem2_22_20, 
        p_wishbone_bd_ram_mem2_22_21, p_wishbone_bd_ram_mem2_22_22, 
        p_wishbone_bd_ram_mem2_22_23, p_wishbone_bd_ram_mem2_23_16, 
        p_wishbone_bd_ram_mem2_23_17, p_wishbone_bd_ram_mem2_23_18, 
        p_wishbone_bd_ram_mem2_23_19, p_wishbone_bd_ram_mem2_23_20, 
        p_wishbone_bd_ram_mem2_23_21, p_wishbone_bd_ram_mem2_23_22, 
        p_wishbone_bd_ram_mem2_23_23, p_wishbone_bd_ram_mem2_24_16, 
        p_wishbone_bd_ram_mem2_24_17, p_wishbone_bd_ram_mem2_24_18, 
        p_wishbone_bd_ram_mem2_24_19, p_wishbone_bd_ram_mem2_24_20, 
        p_wishbone_bd_ram_mem2_24_21, p_wishbone_bd_ram_mem2_24_22, 
        p_wishbone_bd_ram_mem2_24_23, p_wishbone_bd_ram_mem2_25_16, 
        p_wishbone_bd_ram_mem2_25_17, p_wishbone_bd_ram_mem2_25_18, 
        p_wishbone_bd_ram_mem2_25_19, p_wishbone_bd_ram_mem2_25_20, 
        p_wishbone_bd_ram_mem2_25_21, p_wishbone_bd_ram_mem2_25_22, 
        p_wishbone_bd_ram_mem2_25_23, p_wishbone_bd_ram_mem2_26_16, 
        p_wishbone_bd_ram_mem2_26_17, p_wishbone_bd_ram_mem2_26_18, 
        p_wishbone_bd_ram_mem2_26_19, p_wishbone_bd_ram_mem2_26_20, 
        p_wishbone_bd_ram_mem2_26_21, p_wishbone_bd_ram_mem2_26_22, 
        p_wishbone_bd_ram_mem2_26_23, p_wishbone_bd_ram_mem2_27_16, 
        p_wishbone_bd_ram_mem2_27_17, p_wishbone_bd_ram_mem2_27_18, 
        p_wishbone_bd_ram_mem2_27_19, p_wishbone_bd_ram_mem2_27_20, 
        p_wishbone_bd_ram_mem2_27_21, p_wishbone_bd_ram_mem2_27_22, 
        p_wishbone_bd_ram_mem2_27_23, p_wishbone_bd_ram_mem2_28_16, 
        p_wishbone_bd_ram_mem2_28_17, p_wishbone_bd_ram_mem2_28_18, 
        p_wishbone_bd_ram_mem2_28_19, p_wishbone_bd_ram_mem2_28_20, 
        p_wishbone_bd_ram_mem2_28_21, p_wishbone_bd_ram_mem2_28_22, 
        p_wishbone_bd_ram_mem2_28_23, p_wishbone_bd_ram_mem2_29_16, 
        p_wishbone_bd_ram_mem2_29_17, p_wishbone_bd_ram_mem2_29_18, 
        p_wishbone_bd_ram_mem2_29_19, p_wishbone_bd_ram_mem2_29_20, 
        p_wishbone_bd_ram_mem2_29_21, p_wishbone_bd_ram_mem2_29_22, 
        p_wishbone_bd_ram_mem2_29_23, p_wishbone_bd_ram_mem2_30_16, 
        p_wishbone_bd_ram_mem2_30_17, p_wishbone_bd_ram_mem2_30_18, 
        p_wishbone_bd_ram_mem2_30_19, p_wishbone_bd_ram_mem2_30_20, 
        p_wishbone_bd_ram_mem2_30_21, p_wishbone_bd_ram_mem2_30_22, 
        p_wishbone_bd_ram_mem2_30_23, p_wishbone_bd_ram_mem2_31_16, 
        p_wishbone_bd_ram_mem2_31_17, p_wishbone_bd_ram_mem2_31_18, 
        p_wishbone_bd_ram_mem2_31_19, p_wishbone_bd_ram_mem2_31_20, 
        p_wishbone_bd_ram_mem2_31_21, p_wishbone_bd_ram_mem2_31_22, 
        p_wishbone_bd_ram_mem2_31_23, p_wishbone_bd_ram_mem2_32_16, 
        p_wishbone_bd_ram_mem2_32_17, p_wishbone_bd_ram_mem2_32_18, 
        p_wishbone_bd_ram_mem2_32_19, p_wishbone_bd_ram_mem2_32_20, 
        p_wishbone_bd_ram_mem2_32_21, p_wishbone_bd_ram_mem2_32_22, 
        p_wishbone_bd_ram_mem2_32_23, p_wishbone_bd_ram_mem2_33_16, 
        p_wishbone_bd_ram_mem2_33_17, p_wishbone_bd_ram_mem2_33_18, 
        p_wishbone_bd_ram_mem2_33_19, p_wishbone_bd_ram_mem2_33_20, 
        p_wishbone_bd_ram_mem2_33_21, p_wishbone_bd_ram_mem2_33_22, 
        p_wishbone_bd_ram_mem2_33_23, p_wishbone_bd_ram_mem2_34_16, 
        p_wishbone_bd_ram_mem2_34_17, p_wishbone_bd_ram_mem2_34_18, 
        p_wishbone_bd_ram_mem2_34_19, p_wishbone_bd_ram_mem2_34_20, 
        p_wishbone_bd_ram_mem2_34_21, p_wishbone_bd_ram_mem2_34_22, 
        p_wishbone_bd_ram_mem2_34_23, p_wishbone_bd_ram_mem2_35_16, 
        p_wishbone_bd_ram_mem2_35_17, p_wishbone_bd_ram_mem2_35_18, 
        p_wishbone_bd_ram_mem2_35_19, p_wishbone_bd_ram_mem2_35_20, 
        p_wishbone_bd_ram_mem2_35_21, p_wishbone_bd_ram_mem2_35_22, 
        p_wishbone_bd_ram_mem2_35_23, p_wishbone_bd_ram_mem2_36_16, 
        p_wishbone_bd_ram_mem2_36_17, p_wishbone_bd_ram_mem2_36_18, 
        p_wishbone_bd_ram_mem2_36_19, p_wishbone_bd_ram_mem2_36_20, 
        p_wishbone_bd_ram_mem2_36_21, p_wishbone_bd_ram_mem2_36_22, 
        p_wishbone_bd_ram_mem2_36_23, p_wishbone_bd_ram_mem2_37_16, 
        p_wishbone_bd_ram_mem2_37_17, p_wishbone_bd_ram_mem2_37_18, 
        p_wishbone_bd_ram_mem2_37_19, p_wishbone_bd_ram_mem2_37_20, 
        p_wishbone_bd_ram_mem2_37_21, p_wishbone_bd_ram_mem2_37_22, 
        p_wishbone_bd_ram_mem2_37_23, p_wishbone_bd_ram_mem2_38_16, 
        p_wishbone_bd_ram_mem2_38_17, p_wishbone_bd_ram_mem2_38_18, 
        p_wishbone_bd_ram_mem2_38_19, p_wishbone_bd_ram_mem2_38_20, 
        p_wishbone_bd_ram_mem2_38_21, p_wishbone_bd_ram_mem2_38_22, 
        p_wishbone_bd_ram_mem2_38_23, p_wishbone_bd_ram_mem2_39_16, 
        p_wishbone_bd_ram_mem2_39_17, p_wishbone_bd_ram_mem2_39_18, 
        p_wishbone_bd_ram_mem2_39_19, p_wishbone_bd_ram_mem2_39_20, 
        p_wishbone_bd_ram_mem2_39_21, p_wishbone_bd_ram_mem2_39_22, 
        p_wishbone_bd_ram_mem2_39_23, p_wishbone_bd_ram_mem2_40_16, 
        p_wishbone_bd_ram_mem2_40_17, p_wishbone_bd_ram_mem2_40_18, 
        p_wishbone_bd_ram_mem2_40_19, p_wishbone_bd_ram_mem2_40_20, 
        p_wishbone_bd_ram_mem2_40_21, p_wishbone_bd_ram_mem2_40_22, 
        p_wishbone_bd_ram_mem2_40_23, p_wishbone_bd_ram_mem2_41_16, 
        p_wishbone_bd_ram_mem2_41_17, p_wishbone_bd_ram_mem2_41_18, 
        p_wishbone_bd_ram_mem2_41_19, p_wishbone_bd_ram_mem2_41_20, 
        p_wishbone_bd_ram_mem2_41_21, p_wishbone_bd_ram_mem2_41_22, 
        p_wishbone_bd_ram_mem2_41_23, p_wishbone_bd_ram_mem2_42_16, 
        p_wishbone_bd_ram_mem2_42_17, p_wishbone_bd_ram_mem2_42_18, 
        p_wishbone_bd_ram_mem2_42_19, p_wishbone_bd_ram_mem2_42_20, 
        p_wishbone_bd_ram_mem2_42_21, p_wishbone_bd_ram_mem2_42_22, 
        p_wishbone_bd_ram_mem2_42_23, p_wishbone_bd_ram_mem2_43_16, 
        p_wishbone_bd_ram_mem2_43_17, p_wishbone_bd_ram_mem2_43_18, 
        p_wishbone_bd_ram_mem2_43_19, p_wishbone_bd_ram_mem2_43_20, 
        p_wishbone_bd_ram_mem2_43_21, p_wishbone_bd_ram_mem2_43_22, 
        p_wishbone_bd_ram_mem2_43_23, p_wishbone_bd_ram_mem2_44_16, 
        p_wishbone_bd_ram_mem2_44_17, p_wishbone_bd_ram_mem2_44_18, 
        p_wishbone_bd_ram_mem2_44_19, p_wishbone_bd_ram_mem2_44_20, 
        p_wishbone_bd_ram_mem2_44_21, p_wishbone_bd_ram_mem2_44_22, 
        p_wishbone_bd_ram_mem2_44_23, p_wishbone_bd_ram_mem2_45_16, 
        p_wishbone_bd_ram_mem2_45_17, p_wishbone_bd_ram_mem2_45_18, 
        p_wishbone_bd_ram_mem2_45_19, p_wishbone_bd_ram_mem2_45_20, 
        p_wishbone_bd_ram_mem2_45_21, p_wishbone_bd_ram_mem2_45_22, 
        p_wishbone_bd_ram_mem2_45_23, p_wishbone_bd_ram_mem2_46_16, 
        p_wishbone_bd_ram_mem2_46_17, p_wishbone_bd_ram_mem2_46_18, 
        p_wishbone_bd_ram_mem2_46_19, p_wishbone_bd_ram_mem2_46_20, 
        p_wishbone_bd_ram_mem2_46_21, p_wishbone_bd_ram_mem2_46_22, 
        p_wishbone_bd_ram_mem2_46_23, p_wishbone_bd_ram_mem2_47_16, 
        p_wishbone_bd_ram_mem2_47_17, p_wishbone_bd_ram_mem2_47_18, 
        p_wishbone_bd_ram_mem2_47_19, p_wishbone_bd_ram_mem2_47_20, 
        p_wishbone_bd_ram_mem2_47_21, p_wishbone_bd_ram_mem2_47_22, 
        p_wishbone_bd_ram_mem2_47_23, p_wishbone_bd_ram_mem2_48_16, 
        p_wishbone_bd_ram_mem2_48_17, p_wishbone_bd_ram_mem2_48_18, 
        p_wishbone_bd_ram_mem2_48_19, p_wishbone_bd_ram_mem2_48_20, 
        p_wishbone_bd_ram_mem2_48_21, p_wishbone_bd_ram_mem2_48_22, 
        p_wishbone_bd_ram_mem2_48_23, p_wishbone_bd_ram_mem2_49_16, 
        p_wishbone_bd_ram_mem2_49_17, p_wishbone_bd_ram_mem2_49_18, 
        p_wishbone_bd_ram_mem2_49_19, p_wishbone_bd_ram_mem2_49_20, 
        p_wishbone_bd_ram_mem2_49_21, p_wishbone_bd_ram_mem2_49_22, 
        p_wishbone_bd_ram_mem2_49_23, p_wishbone_bd_ram_mem2_50_16, 
        p_wishbone_bd_ram_mem2_50_17, p_wishbone_bd_ram_mem2_50_18, 
        p_wishbone_bd_ram_mem2_50_19, p_wishbone_bd_ram_mem2_50_20, 
        p_wishbone_bd_ram_mem2_50_21, p_wishbone_bd_ram_mem2_50_22, 
        p_wishbone_bd_ram_mem2_50_23, p_wishbone_bd_ram_mem2_51_16, 
        p_wishbone_bd_ram_mem2_51_17, p_wishbone_bd_ram_mem2_51_18, 
        p_wishbone_bd_ram_mem2_51_19, p_wishbone_bd_ram_mem2_51_20, 
        p_wishbone_bd_ram_mem2_51_21, p_wishbone_bd_ram_mem2_51_22, 
        p_wishbone_bd_ram_mem2_51_23, p_wishbone_bd_ram_mem2_52_16, 
        p_wishbone_bd_ram_mem2_52_17, p_wishbone_bd_ram_mem2_52_18, 
        p_wishbone_bd_ram_mem2_52_19, p_wishbone_bd_ram_mem2_52_20, 
        p_wishbone_bd_ram_mem2_52_21, p_wishbone_bd_ram_mem2_52_22, 
        p_wishbone_bd_ram_mem2_52_23, p_wishbone_bd_ram_mem2_53_16, 
        p_wishbone_bd_ram_mem2_53_17, p_wishbone_bd_ram_mem2_53_18, 
        p_wishbone_bd_ram_mem2_53_19, p_wishbone_bd_ram_mem2_53_20, 
        p_wishbone_bd_ram_mem2_53_21, p_wishbone_bd_ram_mem2_53_22, 
        p_wishbone_bd_ram_mem2_53_23, p_wishbone_bd_ram_mem2_54_16, 
        p_wishbone_bd_ram_mem2_54_17, p_wishbone_bd_ram_mem2_54_18, 
        p_wishbone_bd_ram_mem2_54_19, p_wishbone_bd_ram_mem2_54_20, 
        p_wishbone_bd_ram_mem2_54_21, p_wishbone_bd_ram_mem2_54_22, 
        p_wishbone_bd_ram_mem2_54_23, p_wishbone_bd_ram_mem2_55_16, 
        p_wishbone_bd_ram_mem2_55_17, p_wishbone_bd_ram_mem2_55_18, 
        p_wishbone_bd_ram_mem2_55_19, p_wishbone_bd_ram_mem2_55_20, 
        p_wishbone_bd_ram_mem2_55_21, p_wishbone_bd_ram_mem2_55_22, 
        p_wishbone_bd_ram_mem2_55_23, p_wishbone_bd_ram_mem2_56_16, 
        p_wishbone_bd_ram_mem2_56_17, p_wishbone_bd_ram_mem2_56_18, 
        p_wishbone_bd_ram_mem2_56_19, p_wishbone_bd_ram_mem2_56_20, 
        p_wishbone_bd_ram_mem2_56_21, p_wishbone_bd_ram_mem2_56_22, 
        p_wishbone_bd_ram_mem2_56_23, p_wishbone_bd_ram_mem2_57_16, 
        p_wishbone_bd_ram_mem2_57_17, p_wishbone_bd_ram_mem2_57_18, 
        p_wishbone_bd_ram_mem2_57_19, p_wishbone_bd_ram_mem2_57_20, 
        p_wishbone_bd_ram_mem2_57_21, p_wishbone_bd_ram_mem2_57_22, 
        p_wishbone_bd_ram_mem2_57_23, p_wishbone_bd_ram_mem2_58_16, 
        p_wishbone_bd_ram_mem2_58_17, p_wishbone_bd_ram_mem2_58_18, 
        p_wishbone_bd_ram_mem2_58_19, p_wishbone_bd_ram_mem2_58_20, 
        p_wishbone_bd_ram_mem2_58_21, p_wishbone_bd_ram_mem2_58_22, 
        p_wishbone_bd_ram_mem2_58_23, p_wishbone_bd_ram_mem2_59_16, 
        p_wishbone_bd_ram_mem2_59_17, p_wishbone_bd_ram_mem2_59_18, 
        p_wishbone_bd_ram_mem2_59_19, p_wishbone_bd_ram_mem2_59_20, 
        p_wishbone_bd_ram_mem2_59_21, p_wishbone_bd_ram_mem2_59_22, 
        p_wishbone_bd_ram_mem2_59_23, p_wishbone_bd_ram_mem2_60_16, 
        p_wishbone_bd_ram_mem2_60_17, p_wishbone_bd_ram_mem2_60_18, 
        p_wishbone_bd_ram_mem2_60_19, p_wishbone_bd_ram_mem2_60_20, 
        p_wishbone_bd_ram_mem2_60_21, p_wishbone_bd_ram_mem2_60_22, 
        p_wishbone_bd_ram_mem2_60_23, p_wishbone_bd_ram_mem2_61_16, 
        p_wishbone_bd_ram_mem2_61_17, p_wishbone_bd_ram_mem2_61_18, 
        p_wishbone_bd_ram_mem2_61_19, p_wishbone_bd_ram_mem2_61_20, 
        p_wishbone_bd_ram_mem2_61_21, p_wishbone_bd_ram_mem2_61_22, 
        p_wishbone_bd_ram_mem2_61_23, p_wishbone_bd_ram_mem2_62_16, 
        p_wishbone_bd_ram_mem2_62_17, p_wishbone_bd_ram_mem2_62_18, 
        p_wishbone_bd_ram_mem2_62_19, p_wishbone_bd_ram_mem2_62_20, 
        p_wishbone_bd_ram_mem2_62_21, p_wishbone_bd_ram_mem2_62_22, 
        p_wishbone_bd_ram_mem2_62_23, p_wishbone_bd_ram_mem2_63_16, 
        p_wishbone_bd_ram_mem2_63_17, p_wishbone_bd_ram_mem2_63_18, 
        p_wishbone_bd_ram_mem2_63_19, p_wishbone_bd_ram_mem2_63_20, 
        p_wishbone_bd_ram_mem2_63_21, p_wishbone_bd_ram_mem2_63_22, 
        p_wishbone_bd_ram_mem2_63_23, p_wishbone_bd_ram_mem2_64_16, 
        p_wishbone_bd_ram_mem2_64_17, p_wishbone_bd_ram_mem2_64_18, 
        p_wishbone_bd_ram_mem2_64_19, p_wishbone_bd_ram_mem2_64_20, 
        p_wishbone_bd_ram_mem2_64_21, p_wishbone_bd_ram_mem2_64_22, 
        p_wishbone_bd_ram_mem2_64_23, p_wishbone_bd_ram_mem2_65_16, 
        p_wishbone_bd_ram_mem2_65_17, p_wishbone_bd_ram_mem2_65_18, 
        p_wishbone_bd_ram_mem2_65_19, p_wishbone_bd_ram_mem2_65_20, 
        p_wishbone_bd_ram_mem2_65_21, p_wishbone_bd_ram_mem2_65_22, 
        p_wishbone_bd_ram_mem2_65_23, p_wishbone_bd_ram_mem2_66_16, 
        p_wishbone_bd_ram_mem2_66_17, p_wishbone_bd_ram_mem2_66_18, 
        p_wishbone_bd_ram_mem2_66_19, p_wishbone_bd_ram_mem2_66_20, 
        p_wishbone_bd_ram_mem2_66_21, p_wishbone_bd_ram_mem2_66_22, 
        p_wishbone_bd_ram_mem2_66_23, p_wishbone_bd_ram_mem2_67_16, 
        p_wishbone_bd_ram_mem2_67_17, p_wishbone_bd_ram_mem2_67_18, 
        p_wishbone_bd_ram_mem2_67_19, p_wishbone_bd_ram_mem2_67_20, 
        p_wishbone_bd_ram_mem2_67_21, p_wishbone_bd_ram_mem2_67_22, 
        p_wishbone_bd_ram_mem2_67_23, p_wishbone_bd_ram_mem2_68_16, 
        p_wishbone_bd_ram_mem2_68_17, p_wishbone_bd_ram_mem2_68_18, 
        p_wishbone_bd_ram_mem2_68_19, p_wishbone_bd_ram_mem2_68_20, 
        p_wishbone_bd_ram_mem2_68_21, p_wishbone_bd_ram_mem2_68_22, 
        p_wishbone_bd_ram_mem2_68_23, p_wishbone_bd_ram_mem2_69_16, 
        p_wishbone_bd_ram_mem2_69_17, p_wishbone_bd_ram_mem2_69_18, 
        p_wishbone_bd_ram_mem2_69_19, p_wishbone_bd_ram_mem2_69_20, 
        p_wishbone_bd_ram_mem2_69_21, p_wishbone_bd_ram_mem2_69_22, 
        p_wishbone_bd_ram_mem2_69_23, p_wishbone_bd_ram_mem2_70_16, 
        p_wishbone_bd_ram_mem2_70_17, p_wishbone_bd_ram_mem2_70_18, 
        p_wishbone_bd_ram_mem2_70_19, p_wishbone_bd_ram_mem2_70_20, 
        p_wishbone_bd_ram_mem2_70_21, p_wishbone_bd_ram_mem2_70_22, 
        p_wishbone_bd_ram_mem2_70_23, p_wishbone_bd_ram_mem2_71_16, 
        p_wishbone_bd_ram_mem2_71_17, p_wishbone_bd_ram_mem2_71_18, 
        p_wishbone_bd_ram_mem2_71_19, p_wishbone_bd_ram_mem2_71_20, 
        p_wishbone_bd_ram_mem2_71_21, p_wishbone_bd_ram_mem2_71_22, 
        p_wishbone_bd_ram_mem2_71_23, p_wishbone_bd_ram_mem2_72_16, 
        p_wishbone_bd_ram_mem2_72_17, p_wishbone_bd_ram_mem2_72_18, 
        p_wishbone_bd_ram_mem2_72_19, p_wishbone_bd_ram_mem2_72_20, 
        p_wishbone_bd_ram_mem2_72_21, p_wishbone_bd_ram_mem2_72_22, 
        p_wishbone_bd_ram_mem2_72_23, p_wishbone_bd_ram_mem2_73_16, 
        p_wishbone_bd_ram_mem2_73_17, p_wishbone_bd_ram_mem2_73_18, 
        p_wishbone_bd_ram_mem2_73_19, p_wishbone_bd_ram_mem2_73_20, 
        p_wishbone_bd_ram_mem2_73_21, p_wishbone_bd_ram_mem2_73_22, 
        p_wishbone_bd_ram_mem2_73_23, p_wishbone_bd_ram_mem2_74_16, 
        p_wishbone_bd_ram_mem2_74_17, p_wishbone_bd_ram_mem2_74_18, 
        p_wishbone_bd_ram_mem2_74_19, p_wishbone_bd_ram_mem2_74_20, 
        p_wishbone_bd_ram_mem2_74_21, p_wishbone_bd_ram_mem2_74_22, 
        p_wishbone_bd_ram_mem2_74_23, p_wishbone_bd_ram_mem2_75_16, 
        p_wishbone_bd_ram_mem2_75_17, p_wishbone_bd_ram_mem2_75_18, 
        p_wishbone_bd_ram_mem2_75_19, p_wishbone_bd_ram_mem2_75_20, 
        p_wishbone_bd_ram_mem2_75_21, p_wishbone_bd_ram_mem2_75_22, 
        p_wishbone_bd_ram_mem2_75_23, p_wishbone_bd_ram_mem2_76_16, 
        p_wishbone_bd_ram_mem2_76_17, p_wishbone_bd_ram_mem2_76_18, 
        p_wishbone_bd_ram_mem2_76_19, p_wishbone_bd_ram_mem2_76_20, 
        p_wishbone_bd_ram_mem2_76_21, p_wishbone_bd_ram_mem2_76_22, 
        p_wishbone_bd_ram_mem2_76_23, p_wishbone_bd_ram_mem2_77_16, 
        p_wishbone_bd_ram_mem2_77_17, p_wishbone_bd_ram_mem2_77_18, 
        p_wishbone_bd_ram_mem2_77_19, p_wishbone_bd_ram_mem2_77_20, 
        p_wishbone_bd_ram_mem2_77_21, p_wishbone_bd_ram_mem2_77_22, 
        p_wishbone_bd_ram_mem2_77_23, p_wishbone_bd_ram_mem2_78_16, 
        p_wishbone_bd_ram_mem2_78_17, p_wishbone_bd_ram_mem2_78_18, 
        p_wishbone_bd_ram_mem2_78_19, p_wishbone_bd_ram_mem2_78_20, 
        p_wishbone_bd_ram_mem2_78_21, p_wishbone_bd_ram_mem2_78_22, 
        p_wishbone_bd_ram_mem2_78_23, p_wishbone_bd_ram_mem2_79_16, 
        p_wishbone_bd_ram_mem2_79_17, p_wishbone_bd_ram_mem2_79_18, 
        p_wishbone_bd_ram_mem2_79_19, p_wishbone_bd_ram_mem2_79_20, 
        p_wishbone_bd_ram_mem2_79_21, p_wishbone_bd_ram_mem2_79_22, 
        p_wishbone_bd_ram_mem2_79_23, p_wishbone_bd_ram_mem2_80_16, 
        p_wishbone_bd_ram_mem2_80_17, p_wishbone_bd_ram_mem2_80_18, 
        p_wishbone_bd_ram_mem2_80_19, p_wishbone_bd_ram_mem2_80_20, 
        p_wishbone_bd_ram_mem2_80_21, p_wishbone_bd_ram_mem2_80_22, 
        p_wishbone_bd_ram_mem2_80_23, p_wishbone_bd_ram_mem2_81_16, 
        p_wishbone_bd_ram_mem2_81_17, p_wishbone_bd_ram_mem2_81_18, 
        p_wishbone_bd_ram_mem2_81_19, p_wishbone_bd_ram_mem2_81_20, 
        p_wishbone_bd_ram_mem2_81_21, p_wishbone_bd_ram_mem2_81_22, 
        p_wishbone_bd_ram_mem2_81_23, p_wishbone_bd_ram_mem2_82_16, 
        p_wishbone_bd_ram_mem2_82_17, p_wishbone_bd_ram_mem2_82_18, 
        p_wishbone_bd_ram_mem2_82_19, p_wishbone_bd_ram_mem2_82_20, 
        p_wishbone_bd_ram_mem2_82_21, p_wishbone_bd_ram_mem2_82_22, 
        p_wishbone_bd_ram_mem2_82_23, p_wishbone_bd_ram_mem2_83_16, 
        p_wishbone_bd_ram_mem2_83_17, p_wishbone_bd_ram_mem2_83_18, 
        p_wishbone_bd_ram_mem2_83_19, p_wishbone_bd_ram_mem2_83_20, 
        p_wishbone_bd_ram_mem2_83_21, p_wishbone_bd_ram_mem2_83_22, 
        p_wishbone_bd_ram_mem2_83_23, p_wishbone_bd_ram_mem2_84_16, 
        p_wishbone_bd_ram_mem2_84_17, p_wishbone_bd_ram_mem2_84_18, 
        p_wishbone_bd_ram_mem2_84_19, p_wishbone_bd_ram_mem2_84_20, 
        p_wishbone_bd_ram_mem2_84_21, p_wishbone_bd_ram_mem2_84_22, 
        p_wishbone_bd_ram_mem2_84_23, p_wishbone_bd_ram_mem2_85_16, 
        p_wishbone_bd_ram_mem2_85_17, p_wishbone_bd_ram_mem2_85_18, 
        p_wishbone_bd_ram_mem2_85_19, p_wishbone_bd_ram_mem2_85_20, 
        p_wishbone_bd_ram_mem2_85_21, p_wishbone_bd_ram_mem2_85_22, 
        p_wishbone_bd_ram_mem2_85_23, p_wishbone_bd_ram_mem2_86_16, 
        p_wishbone_bd_ram_mem2_86_17, p_wishbone_bd_ram_mem2_86_18, 
        p_wishbone_bd_ram_mem2_86_19, p_wishbone_bd_ram_mem2_86_20, 
        p_wishbone_bd_ram_mem2_86_21, p_wishbone_bd_ram_mem2_86_22, 
        p_wishbone_bd_ram_mem2_86_23, p_wishbone_bd_ram_mem2_87_16, 
        p_wishbone_bd_ram_mem2_87_17, p_wishbone_bd_ram_mem2_87_18, 
        p_wishbone_bd_ram_mem2_87_19, p_wishbone_bd_ram_mem2_87_20, 
        p_wishbone_bd_ram_mem2_87_21, p_wishbone_bd_ram_mem2_87_22, 
        p_wishbone_bd_ram_mem2_87_23, p_wishbone_bd_ram_mem2_88_16, 
        p_wishbone_bd_ram_mem2_88_17, p_wishbone_bd_ram_mem2_88_18, 
        p_wishbone_bd_ram_mem2_88_19, p_wishbone_bd_ram_mem2_88_20, 
        p_wishbone_bd_ram_mem2_88_21, p_wishbone_bd_ram_mem2_88_22, 
        p_wishbone_bd_ram_mem2_88_23, p_wishbone_bd_ram_mem2_89_16, 
        p_wishbone_bd_ram_mem2_89_17, p_wishbone_bd_ram_mem2_89_18, 
        p_wishbone_bd_ram_mem2_89_19, p_wishbone_bd_ram_mem2_89_20, 
        p_wishbone_bd_ram_mem2_89_21, p_wishbone_bd_ram_mem2_89_22, 
        p_wishbone_bd_ram_mem2_89_23, p_wishbone_bd_ram_mem2_90_16, 
        p_wishbone_bd_ram_mem2_90_17, p_wishbone_bd_ram_mem2_90_18, 
        p_wishbone_bd_ram_mem2_90_19, p_wishbone_bd_ram_mem2_90_20, 
        p_wishbone_bd_ram_mem2_90_21, p_wishbone_bd_ram_mem2_90_22, 
        p_wishbone_bd_ram_mem2_90_23, p_wishbone_bd_ram_mem2_91_16, 
        p_wishbone_bd_ram_mem2_91_17, p_wishbone_bd_ram_mem2_91_18, 
        p_wishbone_bd_ram_mem2_91_19, p_wishbone_bd_ram_mem2_91_20, 
        p_wishbone_bd_ram_mem2_91_21, p_wishbone_bd_ram_mem2_91_22, 
        p_wishbone_bd_ram_mem2_91_23, p_wishbone_bd_ram_mem2_92_16, 
        p_wishbone_bd_ram_mem2_92_17, p_wishbone_bd_ram_mem2_92_18, 
        p_wishbone_bd_ram_mem2_92_19, p_wishbone_bd_ram_mem2_92_20, 
        p_wishbone_bd_ram_mem2_92_21, p_wishbone_bd_ram_mem2_92_22, 
        p_wishbone_bd_ram_mem2_92_23, p_wishbone_bd_ram_mem2_93_16, 
        p_wishbone_bd_ram_mem2_93_17, p_wishbone_bd_ram_mem2_93_18, 
        p_wishbone_bd_ram_mem2_93_19, p_wishbone_bd_ram_mem2_93_20, 
        p_wishbone_bd_ram_mem2_93_21, p_wishbone_bd_ram_mem2_93_22, 
        p_wishbone_bd_ram_mem2_93_23, p_wishbone_bd_ram_mem2_94_16, 
        p_wishbone_bd_ram_mem2_94_17, p_wishbone_bd_ram_mem2_94_18, 
        p_wishbone_bd_ram_mem2_94_19, p_wishbone_bd_ram_mem2_94_20, 
        p_wishbone_bd_ram_mem2_94_21, p_wishbone_bd_ram_mem2_94_22, 
        p_wishbone_bd_ram_mem2_94_23, p_wishbone_bd_ram_mem2_95_16, 
        p_wishbone_bd_ram_mem2_95_17, p_wishbone_bd_ram_mem2_95_18, 
        p_wishbone_bd_ram_mem2_95_19, p_wishbone_bd_ram_mem2_95_20, 
        p_wishbone_bd_ram_mem2_95_21, p_wishbone_bd_ram_mem2_95_22, 
        p_wishbone_bd_ram_mem2_95_23, p_wishbone_bd_ram_mem2_96_16, 
        p_wishbone_bd_ram_mem2_96_17, p_wishbone_bd_ram_mem2_96_18, 
        p_wishbone_bd_ram_mem2_96_19, p_wishbone_bd_ram_mem2_96_20, 
        p_wishbone_bd_ram_mem2_96_21, p_wishbone_bd_ram_mem2_96_22, 
        p_wishbone_bd_ram_mem2_96_23, p_wishbone_bd_ram_mem2_97_16, 
        p_wishbone_bd_ram_mem2_97_17, p_wishbone_bd_ram_mem2_97_18, 
        p_wishbone_bd_ram_mem2_97_19, p_wishbone_bd_ram_mem2_97_20, 
        p_wishbone_bd_ram_mem2_97_21, p_wishbone_bd_ram_mem2_97_22, 
        p_wishbone_bd_ram_mem2_97_23, p_wishbone_bd_ram_mem2_98_16, 
        p_wishbone_bd_ram_mem2_98_17, p_wishbone_bd_ram_mem2_98_18, 
        p_wishbone_bd_ram_mem2_98_19, p_wishbone_bd_ram_mem2_98_20, 
        p_wishbone_bd_ram_mem2_98_21, p_wishbone_bd_ram_mem2_98_22, 
        p_wishbone_bd_ram_mem2_98_23, p_wishbone_bd_ram_mem2_99_16, 
        p_wishbone_bd_ram_mem2_99_17, p_wishbone_bd_ram_mem2_99_18, 
        p_wishbone_bd_ram_mem2_99_19, p_wishbone_bd_ram_mem2_99_20, 
        p_wishbone_bd_ram_mem2_99_21, p_wishbone_bd_ram_mem2_99_22, 
        p_wishbone_bd_ram_mem2_99_23, p_wishbone_bd_ram_mem2_100_16, 
        p_wishbone_bd_ram_mem2_100_17, p_wishbone_bd_ram_mem2_100_18, 
        p_wishbone_bd_ram_mem2_100_19, p_wishbone_bd_ram_mem2_100_20, 
        p_wishbone_bd_ram_mem2_100_21, p_wishbone_bd_ram_mem2_100_22, 
        p_wishbone_bd_ram_mem2_100_23, p_wishbone_bd_ram_mem2_101_16, 
        p_wishbone_bd_ram_mem2_101_17, p_wishbone_bd_ram_mem2_101_18, 
        p_wishbone_bd_ram_mem2_101_19, p_wishbone_bd_ram_mem2_101_20, 
        p_wishbone_bd_ram_mem2_101_21, p_wishbone_bd_ram_mem2_101_22, 
        p_wishbone_bd_ram_mem2_101_23, p_wishbone_bd_ram_mem2_102_16, 
        p_wishbone_bd_ram_mem2_102_17, p_wishbone_bd_ram_mem2_102_18, 
        p_wishbone_bd_ram_mem2_102_19, p_wishbone_bd_ram_mem2_102_20, 
        p_wishbone_bd_ram_mem2_102_21, p_wishbone_bd_ram_mem2_102_22, 
        p_wishbone_bd_ram_mem2_102_23, p_wishbone_bd_ram_mem2_103_16, 
        p_wishbone_bd_ram_mem2_103_17, p_wishbone_bd_ram_mem2_103_18, 
        p_wishbone_bd_ram_mem2_103_19, p_wishbone_bd_ram_mem2_103_20, 
        p_wishbone_bd_ram_mem2_103_21, p_wishbone_bd_ram_mem2_103_22, 
        p_wishbone_bd_ram_mem2_103_23, p_wishbone_bd_ram_mem2_104_16, 
        p_wishbone_bd_ram_mem2_104_17, p_wishbone_bd_ram_mem2_104_18, 
        p_wishbone_bd_ram_mem2_104_19, p_wishbone_bd_ram_mem2_104_20, 
        p_wishbone_bd_ram_mem2_104_21, p_wishbone_bd_ram_mem2_104_22, 
        p_wishbone_bd_ram_mem2_104_23, p_wishbone_bd_ram_mem2_105_16, 
        p_wishbone_bd_ram_mem2_105_17, p_wishbone_bd_ram_mem2_105_18, 
        p_wishbone_bd_ram_mem2_105_19, p_wishbone_bd_ram_mem2_105_20, 
        p_wishbone_bd_ram_mem2_105_21, p_wishbone_bd_ram_mem2_105_22, 
        p_wishbone_bd_ram_mem2_105_23, p_wishbone_bd_ram_mem2_106_16, 
        p_wishbone_bd_ram_mem2_106_17, p_wishbone_bd_ram_mem2_106_18, 
        p_wishbone_bd_ram_mem2_106_19, p_wishbone_bd_ram_mem2_106_20, 
        p_wishbone_bd_ram_mem2_106_21, p_wishbone_bd_ram_mem2_106_22, 
        p_wishbone_bd_ram_mem2_106_23, p_wishbone_bd_ram_mem2_107_16, 
        p_wishbone_bd_ram_mem2_107_17, p_wishbone_bd_ram_mem2_107_18, 
        p_wishbone_bd_ram_mem2_107_19, p_wishbone_bd_ram_mem2_107_20, 
        p_wishbone_bd_ram_mem2_107_21, p_wishbone_bd_ram_mem2_107_22, 
        p_wishbone_bd_ram_mem2_107_23, p_wishbone_bd_ram_mem2_108_16, 
        p_wishbone_bd_ram_mem2_108_17, p_wishbone_bd_ram_mem2_108_18, 
        p_wishbone_bd_ram_mem2_108_19, p_wishbone_bd_ram_mem2_108_20, 
        p_wishbone_bd_ram_mem2_108_21, p_wishbone_bd_ram_mem2_108_22, 
        p_wishbone_bd_ram_mem2_108_23, p_wishbone_bd_ram_mem2_109_16, 
        p_wishbone_bd_ram_mem2_109_17, p_wishbone_bd_ram_mem2_109_18, 
        p_wishbone_bd_ram_mem2_109_19, p_wishbone_bd_ram_mem2_109_20, 
        p_wishbone_bd_ram_mem2_109_21, p_wishbone_bd_ram_mem2_109_22, 
        p_wishbone_bd_ram_mem2_109_23, p_wishbone_bd_ram_mem2_110_16, 
        p_wishbone_bd_ram_mem2_110_17, p_wishbone_bd_ram_mem2_110_18, 
        p_wishbone_bd_ram_mem2_110_19, p_wishbone_bd_ram_mem2_110_20, 
        p_wishbone_bd_ram_mem2_110_21, p_wishbone_bd_ram_mem2_110_22, 
        p_wishbone_bd_ram_mem2_110_23, p_wishbone_bd_ram_mem2_111_16, 
        p_wishbone_bd_ram_mem2_111_17, p_wishbone_bd_ram_mem2_111_18, 
        p_wishbone_bd_ram_mem2_111_19, p_wishbone_bd_ram_mem2_111_20, 
        p_wishbone_bd_ram_mem2_111_21, p_wishbone_bd_ram_mem2_111_22, 
        p_wishbone_bd_ram_mem2_111_23, p_wishbone_bd_ram_mem2_112_16, 
        p_wishbone_bd_ram_mem2_112_17, p_wishbone_bd_ram_mem2_112_18, 
        p_wishbone_bd_ram_mem2_112_19, p_wishbone_bd_ram_mem2_112_20, 
        p_wishbone_bd_ram_mem2_112_21, p_wishbone_bd_ram_mem2_112_22, 
        p_wishbone_bd_ram_mem2_112_23, p_wishbone_bd_ram_mem2_113_16, 
        p_wishbone_bd_ram_mem2_113_17, p_wishbone_bd_ram_mem2_113_18, 
        p_wishbone_bd_ram_mem2_113_19, p_wishbone_bd_ram_mem2_113_20, 
        p_wishbone_bd_ram_mem2_113_21, p_wishbone_bd_ram_mem2_113_22, 
        p_wishbone_bd_ram_mem2_113_23, p_wishbone_bd_ram_mem2_114_16, 
        p_wishbone_bd_ram_mem2_114_17, p_wishbone_bd_ram_mem2_114_18, 
        p_wishbone_bd_ram_mem2_114_19, p_wishbone_bd_ram_mem2_114_20, 
        p_wishbone_bd_ram_mem2_114_21, p_wishbone_bd_ram_mem2_114_22, 
        p_wishbone_bd_ram_mem2_114_23, p_wishbone_bd_ram_mem2_115_16, 
        p_wishbone_bd_ram_mem2_115_17, p_wishbone_bd_ram_mem2_115_18, 
        p_wishbone_bd_ram_mem2_115_19, p_wishbone_bd_ram_mem2_115_20, 
        p_wishbone_bd_ram_mem2_115_21, p_wishbone_bd_ram_mem2_115_22, 
        p_wishbone_bd_ram_mem2_115_23, p_wishbone_bd_ram_mem2_116_16, 
        p_wishbone_bd_ram_mem2_116_17, p_wishbone_bd_ram_mem2_116_18, 
        p_wishbone_bd_ram_mem2_116_19, p_wishbone_bd_ram_mem2_116_20, 
        p_wishbone_bd_ram_mem2_116_21, p_wishbone_bd_ram_mem2_116_22, 
        p_wishbone_bd_ram_mem2_116_23, p_wishbone_bd_ram_mem2_117_16, 
        p_wishbone_bd_ram_mem2_117_17, p_wishbone_bd_ram_mem2_117_18, 
        p_wishbone_bd_ram_mem2_117_19, p_wishbone_bd_ram_mem2_117_20, 
        p_wishbone_bd_ram_mem2_117_21, p_wishbone_bd_ram_mem2_117_22, 
        p_wishbone_bd_ram_mem2_117_23, p_wishbone_bd_ram_mem2_118_16, 
        p_wishbone_bd_ram_mem2_118_17, p_wishbone_bd_ram_mem2_118_18, 
        p_wishbone_bd_ram_mem2_118_19, p_wishbone_bd_ram_mem2_118_20, 
        p_wishbone_bd_ram_mem2_118_21, p_wishbone_bd_ram_mem2_118_22, 
        p_wishbone_bd_ram_mem2_118_23, p_wishbone_bd_ram_mem2_119_16, 
        p_wishbone_bd_ram_mem2_119_17, p_wishbone_bd_ram_mem2_119_18, 
        p_wishbone_bd_ram_mem2_119_19, p_wishbone_bd_ram_mem2_119_20, 
        p_wishbone_bd_ram_mem2_119_21, p_wishbone_bd_ram_mem2_119_22, 
        p_wishbone_bd_ram_mem2_119_23, p_wishbone_bd_ram_mem2_120_16, 
        p_wishbone_bd_ram_mem2_120_17, p_wishbone_bd_ram_mem2_120_18, 
        p_wishbone_bd_ram_mem2_120_19, p_wishbone_bd_ram_mem2_120_20, 
        p_wishbone_bd_ram_mem2_120_21, p_wishbone_bd_ram_mem2_120_22, 
        p_wishbone_bd_ram_mem2_120_23, p_wishbone_bd_ram_mem2_121_16, 
        p_wishbone_bd_ram_mem2_121_17, p_wishbone_bd_ram_mem2_121_18, 
        p_wishbone_bd_ram_mem2_121_19, p_wishbone_bd_ram_mem2_121_20, 
        p_wishbone_bd_ram_mem2_121_21, p_wishbone_bd_ram_mem2_121_22, 
        p_wishbone_bd_ram_mem2_121_23, p_wishbone_bd_ram_mem2_122_16, 
        p_wishbone_bd_ram_mem2_122_17, p_wishbone_bd_ram_mem2_122_18, 
        p_wishbone_bd_ram_mem2_122_19, p_wishbone_bd_ram_mem2_122_20, 
        p_wishbone_bd_ram_mem2_122_21, p_wishbone_bd_ram_mem2_122_22, 
        p_wishbone_bd_ram_mem2_122_23, p_wishbone_bd_ram_mem2_123_16, 
        p_wishbone_bd_ram_mem2_123_17, p_wishbone_bd_ram_mem2_123_18, 
        p_wishbone_bd_ram_mem2_123_19, p_wishbone_bd_ram_mem2_123_20, 
        p_wishbone_bd_ram_mem2_123_21, p_wishbone_bd_ram_mem2_123_22, 
        p_wishbone_bd_ram_mem2_123_23, p_wishbone_bd_ram_mem2_124_16, 
        p_wishbone_bd_ram_mem2_124_17, p_wishbone_bd_ram_mem2_124_18, 
        p_wishbone_bd_ram_mem2_124_19, p_wishbone_bd_ram_mem2_124_20, 
        p_wishbone_bd_ram_mem2_124_21, p_wishbone_bd_ram_mem2_124_22, 
        p_wishbone_bd_ram_mem2_124_23, p_wishbone_bd_ram_mem2_125_16, 
        p_wishbone_bd_ram_mem2_125_17, p_wishbone_bd_ram_mem2_125_18, 
        p_wishbone_bd_ram_mem2_125_19, p_wishbone_bd_ram_mem2_125_20, 
        p_wishbone_bd_ram_mem2_125_21, p_wishbone_bd_ram_mem2_125_22, 
        p_wishbone_bd_ram_mem2_125_23, p_wishbone_bd_ram_mem2_126_16, 
        p_wishbone_bd_ram_mem2_126_17, p_wishbone_bd_ram_mem2_126_18, 
        p_wishbone_bd_ram_mem2_126_19, p_wishbone_bd_ram_mem2_126_20, 
        p_wishbone_bd_ram_mem2_126_21, p_wishbone_bd_ram_mem2_126_22, 
        p_wishbone_bd_ram_mem2_126_23, p_wishbone_bd_ram_mem2_127_16, 
        p_wishbone_bd_ram_mem2_127_17, p_wishbone_bd_ram_mem2_127_18, 
        p_wishbone_bd_ram_mem2_127_19, p_wishbone_bd_ram_mem2_127_20, 
        p_wishbone_bd_ram_mem2_127_21, p_wishbone_bd_ram_mem2_127_22, 
        p_wishbone_bd_ram_mem2_127_23, p_wishbone_bd_ram_mem2_128_16, 
        p_wishbone_bd_ram_mem2_128_17, p_wishbone_bd_ram_mem2_128_18, 
        p_wishbone_bd_ram_mem2_128_19, p_wishbone_bd_ram_mem2_128_20, 
        p_wishbone_bd_ram_mem2_128_21, p_wishbone_bd_ram_mem2_128_22, 
        p_wishbone_bd_ram_mem2_128_23, p_wishbone_bd_ram_mem2_129_16, 
        p_wishbone_bd_ram_mem2_129_17, p_wishbone_bd_ram_mem2_129_18, 
        p_wishbone_bd_ram_mem2_129_19, p_wishbone_bd_ram_mem2_129_20, 
        p_wishbone_bd_ram_mem2_129_21, p_wishbone_bd_ram_mem2_129_22, 
        p_wishbone_bd_ram_mem2_129_23, p_wishbone_bd_ram_mem2_130_16, 
        p_wishbone_bd_ram_mem2_130_17, p_wishbone_bd_ram_mem2_130_18, 
        p_wishbone_bd_ram_mem2_130_19, p_wishbone_bd_ram_mem2_130_20, 
        p_wishbone_bd_ram_mem2_130_21, p_wishbone_bd_ram_mem2_130_22, 
        p_wishbone_bd_ram_mem2_130_23, p_wishbone_bd_ram_mem2_131_16, 
        p_wishbone_bd_ram_mem2_131_17, p_wishbone_bd_ram_mem2_131_18, 
        p_wishbone_bd_ram_mem2_131_19, p_wishbone_bd_ram_mem2_131_20, 
        p_wishbone_bd_ram_mem2_131_21, p_wishbone_bd_ram_mem2_131_22, 
        p_wishbone_bd_ram_mem2_131_23, p_wishbone_bd_ram_mem2_132_16, 
        p_wishbone_bd_ram_mem2_132_17, p_wishbone_bd_ram_mem2_132_18, 
        p_wishbone_bd_ram_mem2_132_19, p_wishbone_bd_ram_mem2_132_20, 
        p_wishbone_bd_ram_mem2_132_21, p_wishbone_bd_ram_mem2_132_22, 
        p_wishbone_bd_ram_mem2_132_23, p_wishbone_bd_ram_mem2_133_16, 
        p_wishbone_bd_ram_mem2_133_17, p_wishbone_bd_ram_mem2_133_18, 
        p_wishbone_bd_ram_mem2_133_19, p_wishbone_bd_ram_mem2_133_20, 
        p_wishbone_bd_ram_mem2_133_21, p_wishbone_bd_ram_mem2_133_22, 
        p_wishbone_bd_ram_mem2_133_23, p_wishbone_bd_ram_mem2_134_16, 
        p_wishbone_bd_ram_mem2_134_17, p_wishbone_bd_ram_mem2_134_18, 
        p_wishbone_bd_ram_mem2_134_19, p_wishbone_bd_ram_mem2_134_20, 
        p_wishbone_bd_ram_mem2_134_21, p_wishbone_bd_ram_mem2_134_22, 
        p_wishbone_bd_ram_mem2_134_23, p_wishbone_bd_ram_mem2_135_16, 
        p_wishbone_bd_ram_mem2_135_17, p_wishbone_bd_ram_mem2_135_18, 
        p_wishbone_bd_ram_mem2_135_19, p_wishbone_bd_ram_mem2_135_20, 
        p_wishbone_bd_ram_mem2_135_21, p_wishbone_bd_ram_mem2_135_22, 
        p_wishbone_bd_ram_mem2_135_23, p_wishbone_bd_ram_mem2_136_16, 
        p_wishbone_bd_ram_mem2_136_17, p_wishbone_bd_ram_mem2_136_18, 
        p_wishbone_bd_ram_mem2_136_19, p_wishbone_bd_ram_mem2_136_20, 
        p_wishbone_bd_ram_mem2_136_21, p_wishbone_bd_ram_mem2_136_22, 
        p_wishbone_bd_ram_mem2_136_23, p_wishbone_bd_ram_mem2_137_16, 
        p_wishbone_bd_ram_mem2_137_17, p_wishbone_bd_ram_mem2_137_18, 
        p_wishbone_bd_ram_mem2_137_19, p_wishbone_bd_ram_mem2_137_20, 
        p_wishbone_bd_ram_mem2_137_21, p_wishbone_bd_ram_mem2_137_22, 
        p_wishbone_bd_ram_mem2_137_23, p_wishbone_bd_ram_mem2_138_16, 
        p_wishbone_bd_ram_mem2_138_17, p_wishbone_bd_ram_mem2_138_18, 
        p_wishbone_bd_ram_mem2_138_19, p_wishbone_bd_ram_mem2_138_20, 
        p_wishbone_bd_ram_mem2_138_21, p_wishbone_bd_ram_mem2_138_22, 
        p_wishbone_bd_ram_mem2_138_23, p_wishbone_bd_ram_mem2_139_16, 
        p_wishbone_bd_ram_mem2_139_17, p_wishbone_bd_ram_mem2_139_18, 
        p_wishbone_bd_ram_mem2_139_19, p_wishbone_bd_ram_mem2_139_20, 
        p_wishbone_bd_ram_mem2_139_21, p_wishbone_bd_ram_mem2_139_22, 
        p_wishbone_bd_ram_mem2_139_23, p_wishbone_bd_ram_mem2_140_16, 
        p_wishbone_bd_ram_mem2_140_17, p_wishbone_bd_ram_mem2_140_18, 
        p_wishbone_bd_ram_mem2_140_19, p_wishbone_bd_ram_mem2_140_20, 
        p_wishbone_bd_ram_mem2_140_21, p_wishbone_bd_ram_mem2_140_22, 
        p_wishbone_bd_ram_mem2_140_23, p_wishbone_bd_ram_mem2_141_16, 
        p_wishbone_bd_ram_mem2_141_17, p_wishbone_bd_ram_mem2_141_18, 
        p_wishbone_bd_ram_mem2_141_19, p_wishbone_bd_ram_mem2_141_20, 
        p_wishbone_bd_ram_mem2_141_21, p_wishbone_bd_ram_mem2_141_22, 
        p_wishbone_bd_ram_mem2_141_23, p_wishbone_bd_ram_mem2_142_16, 
        p_wishbone_bd_ram_mem2_142_17, p_wishbone_bd_ram_mem2_142_18, 
        p_wishbone_bd_ram_mem2_142_19, p_wishbone_bd_ram_mem2_142_20, 
        p_wishbone_bd_ram_mem2_142_21, p_wishbone_bd_ram_mem2_142_22, 
        p_wishbone_bd_ram_mem2_142_23, p_wishbone_bd_ram_mem2_143_16, 
        p_wishbone_bd_ram_mem2_143_17, p_wishbone_bd_ram_mem2_143_18, 
        p_wishbone_bd_ram_mem2_143_19, p_wishbone_bd_ram_mem2_143_20, 
        p_wishbone_bd_ram_mem2_143_21, p_wishbone_bd_ram_mem2_143_22, 
        p_wishbone_bd_ram_mem2_143_23, p_wishbone_bd_ram_mem2_144_16, 
        p_wishbone_bd_ram_mem2_144_17, p_wishbone_bd_ram_mem2_144_18, 
        p_wishbone_bd_ram_mem2_144_19, p_wishbone_bd_ram_mem2_144_20, 
        p_wishbone_bd_ram_mem2_144_21, p_wishbone_bd_ram_mem2_144_22, 
        p_wishbone_bd_ram_mem2_144_23, p_wishbone_bd_ram_mem2_145_16, 
        p_wishbone_bd_ram_mem2_145_17, p_wishbone_bd_ram_mem2_145_18, 
        p_wishbone_bd_ram_mem2_145_19, p_wishbone_bd_ram_mem2_145_20, 
        p_wishbone_bd_ram_mem2_145_21, p_wishbone_bd_ram_mem2_145_22, 
        p_wishbone_bd_ram_mem2_145_23, p_wishbone_bd_ram_mem2_146_16, 
        p_wishbone_bd_ram_mem2_146_17, p_wishbone_bd_ram_mem2_146_18, 
        p_wishbone_bd_ram_mem2_146_19, p_wishbone_bd_ram_mem2_146_20, 
        p_wishbone_bd_ram_mem2_146_21, p_wishbone_bd_ram_mem2_146_22, 
        p_wishbone_bd_ram_mem2_146_23, p_wishbone_bd_ram_mem2_147_16, 
        p_wishbone_bd_ram_mem2_147_17, p_wishbone_bd_ram_mem2_147_18, 
        p_wishbone_bd_ram_mem2_147_19, p_wishbone_bd_ram_mem2_147_20, 
        p_wishbone_bd_ram_mem2_147_21, p_wishbone_bd_ram_mem2_147_22, 
        p_wishbone_bd_ram_mem2_147_23, p_wishbone_bd_ram_mem2_148_16, 
        p_wishbone_bd_ram_mem2_148_17, p_wishbone_bd_ram_mem2_148_18, 
        p_wishbone_bd_ram_mem2_148_19, p_wishbone_bd_ram_mem2_148_20, 
        p_wishbone_bd_ram_mem2_148_21, p_wishbone_bd_ram_mem2_148_22, 
        p_wishbone_bd_ram_mem2_148_23, p_wishbone_bd_ram_mem2_149_16, 
        p_wishbone_bd_ram_mem2_149_17, p_wishbone_bd_ram_mem2_149_18, 
        p_wishbone_bd_ram_mem2_149_19, p_wishbone_bd_ram_mem2_149_20, 
        p_wishbone_bd_ram_mem2_149_21, p_wishbone_bd_ram_mem2_149_22, 
        p_wishbone_bd_ram_mem2_149_23, p_wishbone_bd_ram_mem2_150_16, 
        p_wishbone_bd_ram_mem2_150_17, p_wishbone_bd_ram_mem2_150_18, 
        p_wishbone_bd_ram_mem2_150_19, p_wishbone_bd_ram_mem2_150_20, 
        p_wishbone_bd_ram_mem2_150_21, p_wishbone_bd_ram_mem2_150_22, 
        p_wishbone_bd_ram_mem2_150_23, p_wishbone_bd_ram_mem2_151_16, 
        p_wishbone_bd_ram_mem2_151_17, p_wishbone_bd_ram_mem2_151_18, 
        p_wishbone_bd_ram_mem2_151_19, p_wishbone_bd_ram_mem2_151_20, 
        p_wishbone_bd_ram_mem2_151_21, p_wishbone_bd_ram_mem2_151_22, 
        p_wishbone_bd_ram_mem2_151_23, p_wishbone_bd_ram_mem2_152_16, 
        p_wishbone_bd_ram_mem2_152_17, p_wishbone_bd_ram_mem2_152_18, 
        p_wishbone_bd_ram_mem2_152_19, p_wishbone_bd_ram_mem2_152_20, 
        p_wishbone_bd_ram_mem2_152_21, p_wishbone_bd_ram_mem2_152_22, 
        p_wishbone_bd_ram_mem2_152_23, p_wishbone_bd_ram_mem2_153_16, 
        p_wishbone_bd_ram_mem2_153_17, p_wishbone_bd_ram_mem2_153_18, 
        p_wishbone_bd_ram_mem2_153_19, p_wishbone_bd_ram_mem2_153_20, 
        p_wishbone_bd_ram_mem2_153_21, p_wishbone_bd_ram_mem2_153_22, 
        p_wishbone_bd_ram_mem2_153_23, p_wishbone_bd_ram_mem2_154_16, 
        p_wishbone_bd_ram_mem2_154_17, p_wishbone_bd_ram_mem2_154_18, 
        p_wishbone_bd_ram_mem2_154_19, p_wishbone_bd_ram_mem2_154_20, 
        p_wishbone_bd_ram_mem2_154_21, p_wishbone_bd_ram_mem2_154_22, 
        p_wishbone_bd_ram_mem2_154_23, p_wishbone_bd_ram_mem2_155_16, 
        p_wishbone_bd_ram_mem2_155_17, p_wishbone_bd_ram_mem2_155_18, 
        p_wishbone_bd_ram_mem2_155_19, p_wishbone_bd_ram_mem2_155_20, 
        p_wishbone_bd_ram_mem2_155_21, p_wishbone_bd_ram_mem2_155_22, 
        p_wishbone_bd_ram_mem2_155_23, p_wishbone_bd_ram_mem2_156_16, 
        p_wishbone_bd_ram_mem2_156_17, p_wishbone_bd_ram_mem2_156_18, 
        p_wishbone_bd_ram_mem2_156_19, p_wishbone_bd_ram_mem2_156_20, 
        p_wishbone_bd_ram_mem2_156_21, p_wishbone_bd_ram_mem2_156_22, 
        p_wishbone_bd_ram_mem2_156_23, p_wishbone_bd_ram_mem2_157_16, 
        p_wishbone_bd_ram_mem2_157_17, p_wishbone_bd_ram_mem2_157_18, 
        p_wishbone_bd_ram_mem2_157_19, p_wishbone_bd_ram_mem2_157_20, 
        p_wishbone_bd_ram_mem2_157_21, p_wishbone_bd_ram_mem2_157_22, 
        p_wishbone_bd_ram_mem2_157_23, p_wishbone_bd_ram_mem2_158_16, 
        p_wishbone_bd_ram_mem2_158_17, p_wishbone_bd_ram_mem2_158_18, 
        p_wishbone_bd_ram_mem2_158_19, p_wishbone_bd_ram_mem2_158_20, 
        p_wishbone_bd_ram_mem2_158_21, p_wishbone_bd_ram_mem2_158_22, 
        p_wishbone_bd_ram_mem2_158_23, p_wishbone_bd_ram_mem2_159_16, 
        p_wishbone_bd_ram_mem2_159_17, p_wishbone_bd_ram_mem2_159_18, 
        p_wishbone_bd_ram_mem2_159_19, p_wishbone_bd_ram_mem2_159_20, 
        p_wishbone_bd_ram_mem2_159_21, p_wishbone_bd_ram_mem2_159_22, 
        p_wishbone_bd_ram_mem2_159_23, p_wishbone_bd_ram_mem2_160_16, 
        p_wishbone_bd_ram_mem2_160_17, p_wishbone_bd_ram_mem2_160_18, 
        p_wishbone_bd_ram_mem2_160_19, p_wishbone_bd_ram_mem2_160_20, 
        p_wishbone_bd_ram_mem2_160_21, p_wishbone_bd_ram_mem2_160_22, 
        p_wishbone_bd_ram_mem2_160_23, p_wishbone_bd_ram_mem2_161_16, 
        p_wishbone_bd_ram_mem2_161_17, p_wishbone_bd_ram_mem2_161_18, 
        p_wishbone_bd_ram_mem2_161_19, p_wishbone_bd_ram_mem2_161_20, 
        p_wishbone_bd_ram_mem2_161_21, p_wishbone_bd_ram_mem2_161_22, 
        p_wishbone_bd_ram_mem2_161_23, p_wishbone_bd_ram_mem2_162_16, 
        p_wishbone_bd_ram_mem2_162_17, p_wishbone_bd_ram_mem2_162_18, 
        p_wishbone_bd_ram_mem2_162_19, p_wishbone_bd_ram_mem2_162_20, 
        p_wishbone_bd_ram_mem2_162_21, p_wishbone_bd_ram_mem2_162_22, 
        p_wishbone_bd_ram_mem2_162_23, p_wishbone_bd_ram_mem2_163_16, 
        p_wishbone_bd_ram_mem2_163_17, p_wishbone_bd_ram_mem2_163_18, 
        p_wishbone_bd_ram_mem2_163_19, p_wishbone_bd_ram_mem2_163_20, 
        p_wishbone_bd_ram_mem2_163_21, p_wishbone_bd_ram_mem2_163_22, 
        p_wishbone_bd_ram_mem2_163_23, p_wishbone_bd_ram_mem2_164_16, 
        p_wishbone_bd_ram_mem2_164_17, p_wishbone_bd_ram_mem2_164_18, 
        p_wishbone_bd_ram_mem2_164_19, p_wishbone_bd_ram_mem2_164_20, 
        p_wishbone_bd_ram_mem2_164_21, p_wishbone_bd_ram_mem2_164_22, 
        p_wishbone_bd_ram_mem2_164_23, p_wishbone_bd_ram_mem2_165_16, 
        p_wishbone_bd_ram_mem2_165_17, p_wishbone_bd_ram_mem2_165_18, 
        p_wishbone_bd_ram_mem2_165_19, p_wishbone_bd_ram_mem2_165_20, 
        p_wishbone_bd_ram_mem2_165_21, p_wishbone_bd_ram_mem2_165_22, 
        p_wishbone_bd_ram_mem2_165_23, p_wishbone_bd_ram_mem2_166_16, 
        p_wishbone_bd_ram_mem2_166_17, p_wishbone_bd_ram_mem2_166_18, 
        p_wishbone_bd_ram_mem2_166_19, p_wishbone_bd_ram_mem2_166_20, 
        p_wishbone_bd_ram_mem2_166_21, p_wishbone_bd_ram_mem2_166_22, 
        p_wishbone_bd_ram_mem2_166_23, p_wishbone_bd_ram_mem2_167_16, 
        p_wishbone_bd_ram_mem2_167_17, p_wishbone_bd_ram_mem2_167_18, 
        p_wishbone_bd_ram_mem2_167_19, p_wishbone_bd_ram_mem2_167_20, 
        p_wishbone_bd_ram_mem2_167_21, p_wishbone_bd_ram_mem2_167_22, 
        p_wishbone_bd_ram_mem2_167_23, p_wishbone_bd_ram_mem2_168_16, 
        p_wishbone_bd_ram_mem2_168_17, p_wishbone_bd_ram_mem2_168_18, 
        p_wishbone_bd_ram_mem2_168_19, p_wishbone_bd_ram_mem2_168_20, 
        p_wishbone_bd_ram_mem2_168_21, p_wishbone_bd_ram_mem2_168_22, 
        p_wishbone_bd_ram_mem2_168_23, p_wishbone_bd_ram_mem2_169_16, 
        p_wishbone_bd_ram_mem2_169_17, p_wishbone_bd_ram_mem2_169_18, 
        p_wishbone_bd_ram_mem2_169_19, p_wishbone_bd_ram_mem2_169_20, 
        p_wishbone_bd_ram_mem2_169_21, p_wishbone_bd_ram_mem2_169_22, 
        p_wishbone_bd_ram_mem2_169_23, p_wishbone_bd_ram_mem2_170_16, 
        p_wishbone_bd_ram_mem2_170_17, p_wishbone_bd_ram_mem2_170_18, 
        p_wishbone_bd_ram_mem2_170_19, p_wishbone_bd_ram_mem2_170_20, 
        p_wishbone_bd_ram_mem2_170_21, p_wishbone_bd_ram_mem2_170_22, 
        p_wishbone_bd_ram_mem2_170_23, p_wishbone_bd_ram_mem2_171_16, 
        p_wishbone_bd_ram_mem2_171_17, p_wishbone_bd_ram_mem2_171_18, 
        p_wishbone_bd_ram_mem2_171_19, p_wishbone_bd_ram_mem2_171_20, 
        p_wishbone_bd_ram_mem2_171_21, p_wishbone_bd_ram_mem2_171_22, 
        p_wishbone_bd_ram_mem2_171_23, p_wishbone_bd_ram_mem2_172_16, 
        p_wishbone_bd_ram_mem2_172_17, p_wishbone_bd_ram_mem2_172_18, 
        p_wishbone_bd_ram_mem2_172_19, p_wishbone_bd_ram_mem2_172_20, 
        p_wishbone_bd_ram_mem2_172_21, p_wishbone_bd_ram_mem2_172_22, 
        p_wishbone_bd_ram_mem2_172_23, p_wishbone_bd_ram_mem2_173_16, 
        p_wishbone_bd_ram_mem2_173_17, p_wishbone_bd_ram_mem2_173_18, 
        p_wishbone_bd_ram_mem2_173_19, p_wishbone_bd_ram_mem2_173_20, 
        p_wishbone_bd_ram_mem2_173_21, p_wishbone_bd_ram_mem2_173_22, 
        p_wishbone_bd_ram_mem2_173_23, p_wishbone_bd_ram_mem2_174_16, 
        p_wishbone_bd_ram_mem2_174_17, p_wishbone_bd_ram_mem2_174_18, 
        p_wishbone_bd_ram_mem2_174_19, p_wishbone_bd_ram_mem2_174_20, 
        p_wishbone_bd_ram_mem2_174_21, p_wishbone_bd_ram_mem2_174_22, 
        p_wishbone_bd_ram_mem2_174_23, p_wishbone_bd_ram_mem2_175_16, 
        p_wishbone_bd_ram_mem2_175_17, p_wishbone_bd_ram_mem2_175_18, 
        p_wishbone_bd_ram_mem2_175_19, p_wishbone_bd_ram_mem2_175_20, 
        p_wishbone_bd_ram_mem2_175_21, p_wishbone_bd_ram_mem2_175_22, 
        p_wishbone_bd_ram_mem2_175_23, p_wishbone_bd_ram_mem2_176_16, 
        p_wishbone_bd_ram_mem2_176_17, p_wishbone_bd_ram_mem2_176_18, 
        p_wishbone_bd_ram_mem2_176_19, p_wishbone_bd_ram_mem2_176_20, 
        p_wishbone_bd_ram_mem2_176_21, p_wishbone_bd_ram_mem2_176_22, 
        p_wishbone_bd_ram_mem2_176_23, p_wishbone_bd_ram_mem2_177_16, 
        p_wishbone_bd_ram_mem2_177_17, p_wishbone_bd_ram_mem2_177_18, 
        p_wishbone_bd_ram_mem2_177_19, p_wishbone_bd_ram_mem2_177_20, 
        p_wishbone_bd_ram_mem2_177_21, p_wishbone_bd_ram_mem2_177_22, 
        p_wishbone_bd_ram_mem2_177_23, p_wishbone_bd_ram_mem2_178_16, 
        p_wishbone_bd_ram_mem2_178_17, p_wishbone_bd_ram_mem2_178_18, 
        p_wishbone_bd_ram_mem2_178_19, p_wishbone_bd_ram_mem2_178_20, 
        p_wishbone_bd_ram_mem2_178_21, p_wishbone_bd_ram_mem2_178_22, 
        p_wishbone_bd_ram_mem2_178_23, p_wishbone_bd_ram_mem2_179_16, 
        p_wishbone_bd_ram_mem2_179_17, p_wishbone_bd_ram_mem2_179_18, 
        p_wishbone_bd_ram_mem2_179_19, p_wishbone_bd_ram_mem2_179_20, 
        p_wishbone_bd_ram_mem2_179_21, p_wishbone_bd_ram_mem2_179_22, 
        p_wishbone_bd_ram_mem2_179_23, p_wishbone_bd_ram_mem2_180_16, 
        p_wishbone_bd_ram_mem2_180_17, p_wishbone_bd_ram_mem2_180_18, 
        p_wishbone_bd_ram_mem2_180_19, p_wishbone_bd_ram_mem2_180_20, 
        p_wishbone_bd_ram_mem2_180_21, p_wishbone_bd_ram_mem2_180_22, 
        p_wishbone_bd_ram_mem2_180_23, p_wishbone_bd_ram_mem2_181_16, 
        p_wishbone_bd_ram_mem2_181_17, p_wishbone_bd_ram_mem2_181_18, 
        p_wishbone_bd_ram_mem2_181_19, p_wishbone_bd_ram_mem2_181_20, 
        p_wishbone_bd_ram_mem2_181_21, p_wishbone_bd_ram_mem2_181_22, 
        p_wishbone_bd_ram_mem2_181_23, p_wishbone_bd_ram_mem2_182_16, 
        p_wishbone_bd_ram_mem2_182_17, p_wishbone_bd_ram_mem2_182_18, 
        p_wishbone_bd_ram_mem2_182_19, p_wishbone_bd_ram_mem2_182_20, 
        p_wishbone_bd_ram_mem2_182_21, p_wishbone_bd_ram_mem2_182_22, 
        p_wishbone_bd_ram_mem2_182_23, p_wishbone_bd_ram_mem2_183_16, 
        p_wishbone_bd_ram_mem2_183_17, p_wishbone_bd_ram_mem2_183_18, 
        p_wishbone_bd_ram_mem2_183_19, p_wishbone_bd_ram_mem2_183_20, 
        p_wishbone_bd_ram_mem2_183_21, p_wishbone_bd_ram_mem2_183_22, 
        p_wishbone_bd_ram_mem2_183_23, p_wishbone_bd_ram_mem2_184_16, 
        p_wishbone_bd_ram_mem2_184_17, p_wishbone_bd_ram_mem2_184_18, 
        p_wishbone_bd_ram_mem2_184_19, p_wishbone_bd_ram_mem2_184_20, 
        p_wishbone_bd_ram_mem2_184_21, p_wishbone_bd_ram_mem2_184_22, 
        p_wishbone_bd_ram_mem2_184_23, p_wishbone_bd_ram_mem2_185_16, 
        p_wishbone_bd_ram_mem2_185_17, p_wishbone_bd_ram_mem2_185_18, 
        p_wishbone_bd_ram_mem2_185_19, p_wishbone_bd_ram_mem2_185_20, 
        p_wishbone_bd_ram_mem2_185_21, p_wishbone_bd_ram_mem2_185_22, 
        p_wishbone_bd_ram_mem2_185_23, p_wishbone_bd_ram_mem2_186_16, 
        p_wishbone_bd_ram_mem2_186_17, p_wishbone_bd_ram_mem2_186_18, 
        p_wishbone_bd_ram_mem2_186_19, p_wishbone_bd_ram_mem2_186_20, 
        p_wishbone_bd_ram_mem2_186_21, p_wishbone_bd_ram_mem2_186_22, 
        p_wishbone_bd_ram_mem2_186_23, p_wishbone_bd_ram_mem2_187_16, 
        p_wishbone_bd_ram_mem2_187_17, p_wishbone_bd_ram_mem2_187_18, 
        p_wishbone_bd_ram_mem2_187_19, p_wishbone_bd_ram_mem2_187_20, 
        p_wishbone_bd_ram_mem2_187_21, p_wishbone_bd_ram_mem2_187_22, 
        p_wishbone_bd_ram_mem2_187_23, p_wishbone_bd_ram_mem2_188_16, 
        p_wishbone_bd_ram_mem2_188_17, p_wishbone_bd_ram_mem2_188_18, 
        p_wishbone_bd_ram_mem2_188_19, p_wishbone_bd_ram_mem2_188_20, 
        p_wishbone_bd_ram_mem2_188_21, p_wishbone_bd_ram_mem2_188_22, 
        p_wishbone_bd_ram_mem2_188_23, p_wishbone_bd_ram_mem2_189_16, 
        p_wishbone_bd_ram_mem2_189_17, p_wishbone_bd_ram_mem2_189_18, 
        p_wishbone_bd_ram_mem2_189_19, p_wishbone_bd_ram_mem2_189_20, 
        p_wishbone_bd_ram_mem2_189_21, p_wishbone_bd_ram_mem2_189_22, 
        p_wishbone_bd_ram_mem2_189_23, p_wishbone_bd_ram_mem2_190_16, 
        p_wishbone_bd_ram_mem2_190_17, p_wishbone_bd_ram_mem2_190_18, 
        p_wishbone_bd_ram_mem2_190_19, p_wishbone_bd_ram_mem2_190_20, 
        p_wishbone_bd_ram_mem2_190_21, p_wishbone_bd_ram_mem2_190_22, 
        p_wishbone_bd_ram_mem2_190_23, p_wishbone_bd_ram_mem2_191_16, 
        p_wishbone_bd_ram_mem2_191_17, p_wishbone_bd_ram_mem2_191_18, 
        p_wishbone_bd_ram_mem2_191_19, p_wishbone_bd_ram_mem2_191_20, 
        p_wishbone_bd_ram_mem2_191_21, p_wishbone_bd_ram_mem2_191_22, 
        p_wishbone_bd_ram_mem2_191_23, p_wishbone_bd_ram_mem2_192_16, 
        p_wishbone_bd_ram_mem2_192_17, p_wishbone_bd_ram_mem2_192_18, 
        p_wishbone_bd_ram_mem2_192_19, p_wishbone_bd_ram_mem2_192_20, 
        p_wishbone_bd_ram_mem2_192_21, p_wishbone_bd_ram_mem2_192_22, 
        p_wishbone_bd_ram_mem2_192_23, p_wishbone_bd_ram_mem2_193_16, 
        p_wishbone_bd_ram_mem2_193_17, p_wishbone_bd_ram_mem2_193_18, 
        p_wishbone_bd_ram_mem2_193_19, p_wishbone_bd_ram_mem2_193_20, 
        p_wishbone_bd_ram_mem2_193_21, p_wishbone_bd_ram_mem2_193_22, 
        p_wishbone_bd_ram_mem2_193_23, p_wishbone_bd_ram_mem2_194_16, 
        p_wishbone_bd_ram_mem2_194_17, p_wishbone_bd_ram_mem2_194_18, 
        p_wishbone_bd_ram_mem2_194_19, p_wishbone_bd_ram_mem2_194_20, 
        p_wishbone_bd_ram_mem2_194_21, p_wishbone_bd_ram_mem2_194_22, 
        p_wishbone_bd_ram_mem2_194_23, p_wishbone_bd_ram_mem2_195_16, 
        p_wishbone_bd_ram_mem2_195_17, p_wishbone_bd_ram_mem2_195_18, 
        p_wishbone_bd_ram_mem2_195_19, p_wishbone_bd_ram_mem2_195_20, 
        p_wishbone_bd_ram_mem2_195_21, p_wishbone_bd_ram_mem2_195_22, 
        p_wishbone_bd_ram_mem2_195_23, p_wishbone_bd_ram_mem2_196_16, 
        p_wishbone_bd_ram_mem2_196_17, p_wishbone_bd_ram_mem2_196_18, 
        p_wishbone_bd_ram_mem2_196_19, p_wishbone_bd_ram_mem2_196_20, 
        p_wishbone_bd_ram_mem2_196_21, p_wishbone_bd_ram_mem2_196_22, 
        p_wishbone_bd_ram_mem2_196_23, p_wishbone_bd_ram_mem2_197_16, 
        p_wishbone_bd_ram_mem2_197_17, p_wishbone_bd_ram_mem2_197_18, 
        p_wishbone_bd_ram_mem2_197_19, p_wishbone_bd_ram_mem2_197_20, 
        p_wishbone_bd_ram_mem2_197_21, p_wishbone_bd_ram_mem2_197_22, 
        p_wishbone_bd_ram_mem2_197_23, p_wishbone_bd_ram_mem2_198_16, 
        p_wishbone_bd_ram_mem2_198_17, p_wishbone_bd_ram_mem2_198_18, 
        p_wishbone_bd_ram_mem2_198_19, p_wishbone_bd_ram_mem2_198_20, 
        p_wishbone_bd_ram_mem2_198_21, p_wishbone_bd_ram_mem2_198_22, 
        p_wishbone_bd_ram_mem2_198_23, p_wishbone_bd_ram_mem2_199_16, 
        p_wishbone_bd_ram_mem2_199_17, p_wishbone_bd_ram_mem2_199_18, 
        p_wishbone_bd_ram_mem2_199_19, p_wishbone_bd_ram_mem2_199_20, 
        p_wishbone_bd_ram_mem2_199_21, p_wishbone_bd_ram_mem2_199_22, 
        p_wishbone_bd_ram_mem2_199_23, p_wishbone_bd_ram_mem2_200_16, 
        p_wishbone_bd_ram_mem2_200_17, p_wishbone_bd_ram_mem2_200_18, 
        p_wishbone_bd_ram_mem2_200_19, p_wishbone_bd_ram_mem2_200_20, 
        p_wishbone_bd_ram_mem2_200_21, p_wishbone_bd_ram_mem2_200_22, 
        p_wishbone_bd_ram_mem2_200_23, p_wishbone_bd_ram_mem2_201_16, 
        p_wishbone_bd_ram_mem2_201_17, p_wishbone_bd_ram_mem2_201_18, 
        p_wishbone_bd_ram_mem2_201_19, p_wishbone_bd_ram_mem2_201_20, 
        p_wishbone_bd_ram_mem2_201_21, p_wishbone_bd_ram_mem2_201_22, 
        p_wishbone_bd_ram_mem2_201_23, p_wishbone_bd_ram_mem2_202_16, 
        p_wishbone_bd_ram_mem2_202_17, p_wishbone_bd_ram_mem2_202_18, 
        p_wishbone_bd_ram_mem2_202_19, p_wishbone_bd_ram_mem2_202_20, 
        p_wishbone_bd_ram_mem2_202_21, p_wishbone_bd_ram_mem2_202_22, 
        p_wishbone_bd_ram_mem2_202_23, p_wishbone_bd_ram_mem2_203_16, 
        p_wishbone_bd_ram_mem2_203_17, p_wishbone_bd_ram_mem2_203_18, 
        p_wishbone_bd_ram_mem2_203_19, p_wishbone_bd_ram_mem2_203_20, 
        p_wishbone_bd_ram_mem2_203_21, p_wishbone_bd_ram_mem2_203_22, 
        p_wishbone_bd_ram_mem2_203_23, p_wishbone_bd_ram_mem2_204_16, 
        p_wishbone_bd_ram_mem2_204_17, p_wishbone_bd_ram_mem2_204_18, 
        p_wishbone_bd_ram_mem2_204_19, p_wishbone_bd_ram_mem2_204_20, 
        p_wishbone_bd_ram_mem2_204_21, p_wishbone_bd_ram_mem2_204_22, 
        p_wishbone_bd_ram_mem2_204_23, p_wishbone_bd_ram_mem2_205_16, 
        p_wishbone_bd_ram_mem2_205_17, p_wishbone_bd_ram_mem2_205_18, 
        p_wishbone_bd_ram_mem2_205_19, p_wishbone_bd_ram_mem2_205_20, 
        p_wishbone_bd_ram_mem2_205_21, p_wishbone_bd_ram_mem2_205_22, 
        p_wishbone_bd_ram_mem2_205_23, p_wishbone_bd_ram_mem2_206_16, 
        p_wishbone_bd_ram_mem2_206_17, p_wishbone_bd_ram_mem2_206_18, 
        p_wishbone_bd_ram_mem2_206_19, p_wishbone_bd_ram_mem2_206_20, 
        p_wishbone_bd_ram_mem2_206_21, p_wishbone_bd_ram_mem2_206_22, 
        p_wishbone_bd_ram_mem2_206_23, p_wishbone_bd_ram_mem2_207_16, 
        p_wishbone_bd_ram_mem2_207_17, p_wishbone_bd_ram_mem2_207_18, 
        p_wishbone_bd_ram_mem2_207_19, p_wishbone_bd_ram_mem2_207_20, 
        p_wishbone_bd_ram_mem2_207_21, p_wishbone_bd_ram_mem2_207_22, 
        p_wishbone_bd_ram_mem2_207_23, p_wishbone_bd_ram_mem2_208_16, 
        p_wishbone_bd_ram_mem2_208_17, p_wishbone_bd_ram_mem2_208_18, 
        p_wishbone_bd_ram_mem2_208_19, p_wishbone_bd_ram_mem2_208_20, 
        p_wishbone_bd_ram_mem2_208_21, p_wishbone_bd_ram_mem2_208_22, 
        p_wishbone_bd_ram_mem2_208_23, p_wishbone_bd_ram_mem2_209_16, 
        p_wishbone_bd_ram_mem2_209_17, p_wishbone_bd_ram_mem2_209_18, 
        p_wishbone_bd_ram_mem2_209_19, p_wishbone_bd_ram_mem2_209_20, 
        p_wishbone_bd_ram_mem2_209_21, p_wishbone_bd_ram_mem2_209_22, 
        p_wishbone_bd_ram_mem2_209_23, p_wishbone_bd_ram_mem2_210_16, 
        p_wishbone_bd_ram_mem2_210_17, p_wishbone_bd_ram_mem2_210_18, 
        p_wishbone_bd_ram_mem2_210_19, p_wishbone_bd_ram_mem2_210_20, 
        p_wishbone_bd_ram_mem2_210_21, p_wishbone_bd_ram_mem2_210_22, 
        p_wishbone_bd_ram_mem2_210_23, p_wishbone_bd_ram_mem2_211_16, 
        p_wishbone_bd_ram_mem2_211_17, p_wishbone_bd_ram_mem2_211_18, 
        p_wishbone_bd_ram_mem2_211_19, p_wishbone_bd_ram_mem2_211_20, 
        p_wishbone_bd_ram_mem2_211_21, p_wishbone_bd_ram_mem2_211_22, 
        p_wishbone_bd_ram_mem2_211_23, p_wishbone_bd_ram_mem2_212_16, 
        p_wishbone_bd_ram_mem2_212_17, p_wishbone_bd_ram_mem2_212_18, 
        p_wishbone_bd_ram_mem2_212_19, p_wishbone_bd_ram_mem2_212_20, 
        p_wishbone_bd_ram_mem2_212_21, p_wishbone_bd_ram_mem2_212_22, 
        p_wishbone_bd_ram_mem2_212_23, p_wishbone_bd_ram_mem2_213_16, 
        p_wishbone_bd_ram_mem2_213_17, p_wishbone_bd_ram_mem2_213_18, 
        p_wishbone_bd_ram_mem2_213_19, p_wishbone_bd_ram_mem2_213_20, 
        p_wishbone_bd_ram_mem2_213_21, p_wishbone_bd_ram_mem2_213_22, 
        p_wishbone_bd_ram_mem2_213_23, p_wishbone_bd_ram_mem2_214_16, 
        p_wishbone_bd_ram_mem2_214_17, p_wishbone_bd_ram_mem2_214_18, 
        p_wishbone_bd_ram_mem2_214_19, p_wishbone_bd_ram_mem2_214_20, 
        p_wishbone_bd_ram_mem2_214_21, p_wishbone_bd_ram_mem2_214_22, 
        p_wishbone_bd_ram_mem2_214_23, p_wishbone_bd_ram_mem2_215_16, 
        p_wishbone_bd_ram_mem2_215_17, p_wishbone_bd_ram_mem2_215_18, 
        p_wishbone_bd_ram_mem2_215_19, p_wishbone_bd_ram_mem2_215_20, 
        p_wishbone_bd_ram_mem2_215_21, p_wishbone_bd_ram_mem2_215_22, 
        p_wishbone_bd_ram_mem2_215_23, p_wishbone_bd_ram_mem2_216_16, 
        p_wishbone_bd_ram_mem2_216_17, p_wishbone_bd_ram_mem2_216_18, 
        p_wishbone_bd_ram_mem2_216_19, p_wishbone_bd_ram_mem2_216_20, 
        p_wishbone_bd_ram_mem2_216_21, p_wishbone_bd_ram_mem2_216_22, 
        p_wishbone_bd_ram_mem2_216_23, p_wishbone_bd_ram_mem2_217_16, 
        p_wishbone_bd_ram_mem2_217_17, p_wishbone_bd_ram_mem2_217_18, 
        p_wishbone_bd_ram_mem2_217_19, p_wishbone_bd_ram_mem2_217_20, 
        p_wishbone_bd_ram_mem2_217_21, p_wishbone_bd_ram_mem2_217_22, 
        p_wishbone_bd_ram_mem2_217_23, p_wishbone_bd_ram_mem2_218_16, 
        p_wishbone_bd_ram_mem2_218_17, p_wishbone_bd_ram_mem2_218_18, 
        p_wishbone_bd_ram_mem2_218_19, p_wishbone_bd_ram_mem2_218_20, 
        p_wishbone_bd_ram_mem2_218_21, p_wishbone_bd_ram_mem2_218_22, 
        p_wishbone_bd_ram_mem2_218_23, p_wishbone_bd_ram_mem2_219_16, 
        p_wishbone_bd_ram_mem2_219_17, p_wishbone_bd_ram_mem2_219_18, 
        p_wishbone_bd_ram_mem2_219_19, p_wishbone_bd_ram_mem2_219_20, 
        p_wishbone_bd_ram_mem2_219_21, p_wishbone_bd_ram_mem2_219_22, 
        p_wishbone_bd_ram_mem2_219_23, p_wishbone_bd_ram_mem2_220_16, 
        p_wishbone_bd_ram_mem2_220_17, p_wishbone_bd_ram_mem2_220_18, 
        p_wishbone_bd_ram_mem2_220_19, p_wishbone_bd_ram_mem2_220_20, 
        p_wishbone_bd_ram_mem2_220_21, p_wishbone_bd_ram_mem2_220_22, 
        p_wishbone_bd_ram_mem2_220_23, p_wishbone_bd_ram_mem2_221_16, 
        p_wishbone_bd_ram_mem2_221_17, p_wishbone_bd_ram_mem2_221_18, 
        p_wishbone_bd_ram_mem2_221_19, p_wishbone_bd_ram_mem2_221_20, 
        p_wishbone_bd_ram_mem2_221_21, p_wishbone_bd_ram_mem2_221_22, 
        p_wishbone_bd_ram_mem2_221_23, p_wishbone_bd_ram_mem2_222_16, 
        p_wishbone_bd_ram_mem2_222_17, p_wishbone_bd_ram_mem2_222_18, 
        p_wishbone_bd_ram_mem2_222_19, p_wishbone_bd_ram_mem2_222_20, 
        p_wishbone_bd_ram_mem2_222_21, p_wishbone_bd_ram_mem2_222_22, 
        p_wishbone_bd_ram_mem2_222_23, p_wishbone_bd_ram_mem2_223_16, 
        p_wishbone_bd_ram_mem2_223_17, p_wishbone_bd_ram_mem2_223_18, 
        p_wishbone_bd_ram_mem2_223_19, p_wishbone_bd_ram_mem2_223_20, 
        p_wishbone_bd_ram_mem2_223_21, p_wishbone_bd_ram_mem2_223_22, 
        p_wishbone_bd_ram_mem2_223_23, p_wishbone_bd_ram_mem2_224_16, 
        p_wishbone_bd_ram_mem2_224_17, p_wishbone_bd_ram_mem2_224_18, 
        p_wishbone_bd_ram_mem2_224_19, p_wishbone_bd_ram_mem2_224_20, 
        p_wishbone_bd_ram_mem2_224_21, p_wishbone_bd_ram_mem2_224_22, 
        p_wishbone_bd_ram_mem2_224_23, p_wishbone_bd_ram_mem2_225_16, 
        p_wishbone_bd_ram_mem2_225_17, p_wishbone_bd_ram_mem2_225_18, 
        p_wishbone_bd_ram_mem2_225_19, p_wishbone_bd_ram_mem2_225_20, 
        p_wishbone_bd_ram_mem2_225_21, p_wishbone_bd_ram_mem2_225_22, 
        p_wishbone_bd_ram_mem2_225_23, p_wishbone_bd_ram_mem2_226_16, 
        p_wishbone_bd_ram_mem2_226_17, p_wishbone_bd_ram_mem2_226_18, 
        p_wishbone_bd_ram_mem2_226_19, p_wishbone_bd_ram_mem2_226_20, 
        p_wishbone_bd_ram_mem2_226_21, p_wishbone_bd_ram_mem2_226_22, 
        p_wishbone_bd_ram_mem2_226_23, p_wishbone_bd_ram_mem2_227_16, 
        p_wishbone_bd_ram_mem2_227_17, p_wishbone_bd_ram_mem2_227_18, 
        p_wishbone_bd_ram_mem2_227_19, p_wishbone_bd_ram_mem2_227_20, 
        p_wishbone_bd_ram_mem2_227_21, p_wishbone_bd_ram_mem2_227_22, 
        p_wishbone_bd_ram_mem2_227_23, p_wishbone_bd_ram_mem2_228_16, 
        p_wishbone_bd_ram_mem2_228_17, p_wishbone_bd_ram_mem2_228_18, 
        p_wishbone_bd_ram_mem2_228_19, p_wishbone_bd_ram_mem2_228_20, 
        p_wishbone_bd_ram_mem2_228_21, p_wishbone_bd_ram_mem2_228_22, 
        p_wishbone_bd_ram_mem2_228_23, p_wishbone_bd_ram_mem2_229_16, 
        p_wishbone_bd_ram_mem2_229_17, p_wishbone_bd_ram_mem2_229_18, 
        p_wishbone_bd_ram_mem2_229_19, p_wishbone_bd_ram_mem2_229_20, 
        p_wishbone_bd_ram_mem2_229_21, p_wishbone_bd_ram_mem2_229_22, 
        p_wishbone_bd_ram_mem2_229_23, p_wishbone_bd_ram_mem2_230_16, 
        p_wishbone_bd_ram_mem2_230_17, p_wishbone_bd_ram_mem2_230_18, 
        p_wishbone_bd_ram_mem2_230_19, p_wishbone_bd_ram_mem2_230_20, 
        p_wishbone_bd_ram_mem2_230_21, p_wishbone_bd_ram_mem2_230_22, 
        p_wishbone_bd_ram_mem2_230_23, p_wishbone_bd_ram_mem2_231_16, 
        p_wishbone_bd_ram_mem2_231_17, p_wishbone_bd_ram_mem2_231_18, 
        p_wishbone_bd_ram_mem2_231_19, p_wishbone_bd_ram_mem2_231_20, 
        p_wishbone_bd_ram_mem2_231_21, p_wishbone_bd_ram_mem2_231_22, 
        p_wishbone_bd_ram_mem2_231_23, p_wishbone_bd_ram_mem2_232_16, 
        p_wishbone_bd_ram_mem2_232_17, p_wishbone_bd_ram_mem2_232_18, 
        p_wishbone_bd_ram_mem2_232_19, p_wishbone_bd_ram_mem2_232_20, 
        p_wishbone_bd_ram_mem2_232_21, p_wishbone_bd_ram_mem2_232_22, 
        p_wishbone_bd_ram_mem2_232_23, p_wishbone_bd_ram_mem2_233_16, 
        p_wishbone_bd_ram_mem2_233_17, p_wishbone_bd_ram_mem2_233_18, 
        p_wishbone_bd_ram_mem2_233_19, p_wishbone_bd_ram_mem2_233_20, 
        p_wishbone_bd_ram_mem2_233_21, p_wishbone_bd_ram_mem2_233_22, 
        p_wishbone_bd_ram_mem2_233_23, p_wishbone_bd_ram_mem2_234_16, 
        p_wishbone_bd_ram_mem2_234_17, p_wishbone_bd_ram_mem2_234_18, 
        p_wishbone_bd_ram_mem2_234_19, p_wishbone_bd_ram_mem2_234_20, 
        p_wishbone_bd_ram_mem2_234_21, p_wishbone_bd_ram_mem2_234_22, 
        p_wishbone_bd_ram_mem2_234_23, p_wishbone_bd_ram_mem2_235_16, 
        p_wishbone_bd_ram_mem2_235_17, p_wishbone_bd_ram_mem2_235_18, 
        p_wishbone_bd_ram_mem2_235_19, p_wishbone_bd_ram_mem2_235_20, 
        p_wishbone_bd_ram_mem2_235_21, p_wishbone_bd_ram_mem2_235_22, 
        p_wishbone_bd_ram_mem2_235_23, p_wishbone_bd_ram_mem2_236_16, 
        p_wishbone_bd_ram_mem2_236_17, p_wishbone_bd_ram_mem2_236_18, 
        p_wishbone_bd_ram_mem2_236_19, p_wishbone_bd_ram_mem2_236_20, 
        p_wishbone_bd_ram_mem2_236_21, p_wishbone_bd_ram_mem2_236_22, 
        p_wishbone_bd_ram_mem2_236_23, p_wishbone_bd_ram_mem2_237_16, 
        p_wishbone_bd_ram_mem2_237_17, p_wishbone_bd_ram_mem2_237_18, 
        p_wishbone_bd_ram_mem2_237_19, p_wishbone_bd_ram_mem2_237_20, 
        p_wishbone_bd_ram_mem2_237_21, p_wishbone_bd_ram_mem2_237_22, 
        p_wishbone_bd_ram_mem2_237_23, p_wishbone_bd_ram_mem2_238_16, 
        p_wishbone_bd_ram_mem2_238_17, p_wishbone_bd_ram_mem2_238_18, 
        p_wishbone_bd_ram_mem2_238_19, p_wishbone_bd_ram_mem2_238_20, 
        p_wishbone_bd_ram_mem2_238_21, p_wishbone_bd_ram_mem2_238_22, 
        p_wishbone_bd_ram_mem2_238_23, p_wishbone_bd_ram_mem2_239_16, 
        p_wishbone_bd_ram_mem2_239_17, p_wishbone_bd_ram_mem2_239_18, 
        p_wishbone_bd_ram_mem2_239_19, p_wishbone_bd_ram_mem2_239_20, 
        p_wishbone_bd_ram_mem2_239_21, p_wishbone_bd_ram_mem2_239_22, 
        p_wishbone_bd_ram_mem2_239_23, p_wishbone_bd_ram_mem2_240_16, 
        p_wishbone_bd_ram_mem2_240_17, p_wishbone_bd_ram_mem2_240_18, 
        p_wishbone_bd_ram_mem2_240_19, p_wishbone_bd_ram_mem2_240_20, 
        p_wishbone_bd_ram_mem2_240_21, p_wishbone_bd_ram_mem2_240_22, 
        p_wishbone_bd_ram_mem2_240_23, p_wishbone_bd_ram_mem2_241_16, 
        p_wishbone_bd_ram_mem2_241_17, p_wishbone_bd_ram_mem2_241_18, 
        p_wishbone_bd_ram_mem2_241_19, p_wishbone_bd_ram_mem2_241_20, 
        p_wishbone_bd_ram_mem2_241_21, p_wishbone_bd_ram_mem2_241_22, 
        p_wishbone_bd_ram_mem2_241_23, p_wishbone_bd_ram_mem2_242_16, 
        p_wishbone_bd_ram_mem2_242_17, p_wishbone_bd_ram_mem2_242_18, 
        p_wishbone_bd_ram_mem2_242_19, p_wishbone_bd_ram_mem2_242_20, 
        p_wishbone_bd_ram_mem2_242_21, p_wishbone_bd_ram_mem2_242_22, 
        p_wishbone_bd_ram_mem2_242_23, p_wishbone_bd_ram_mem2_243_16, 
        p_wishbone_bd_ram_mem2_243_17, p_wishbone_bd_ram_mem2_243_18, 
        p_wishbone_bd_ram_mem2_243_19, p_wishbone_bd_ram_mem2_243_20, 
        p_wishbone_bd_ram_mem2_243_21, p_wishbone_bd_ram_mem2_243_22, 
        p_wishbone_bd_ram_mem2_243_23, p_wishbone_bd_ram_mem2_244_16, 
        p_wishbone_bd_ram_mem2_244_17, p_wishbone_bd_ram_mem2_244_18, 
        p_wishbone_bd_ram_mem2_244_19, p_wishbone_bd_ram_mem2_244_20, 
        p_wishbone_bd_ram_mem2_244_21, p_wishbone_bd_ram_mem2_244_22, 
        p_wishbone_bd_ram_mem2_244_23, p_wishbone_bd_ram_mem2_245_16, 
        p_wishbone_bd_ram_mem2_245_17, p_wishbone_bd_ram_mem2_245_18, 
        p_wishbone_bd_ram_mem2_245_19, p_wishbone_bd_ram_mem2_245_20, 
        p_wishbone_bd_ram_mem2_245_21, p_wishbone_bd_ram_mem2_245_22, 
        p_wishbone_bd_ram_mem2_245_23, p_wishbone_bd_ram_mem2_246_16, 
        p_wishbone_bd_ram_mem2_246_17, p_wishbone_bd_ram_mem2_246_18, 
        p_wishbone_bd_ram_mem2_246_19, p_wishbone_bd_ram_mem2_246_20, 
        p_wishbone_bd_ram_mem2_246_21, p_wishbone_bd_ram_mem2_246_22, 
        p_wishbone_bd_ram_mem2_246_23, p_wishbone_bd_ram_mem2_247_16, 
        p_wishbone_bd_ram_mem2_247_17, p_wishbone_bd_ram_mem2_247_18, 
        p_wishbone_bd_ram_mem2_247_19, p_wishbone_bd_ram_mem2_247_20, 
        p_wishbone_bd_ram_mem2_247_21, p_wishbone_bd_ram_mem2_247_22, 
        p_wishbone_bd_ram_mem2_247_23, p_wishbone_bd_ram_mem2_248_16, 
        p_wishbone_bd_ram_mem2_248_17, p_wishbone_bd_ram_mem2_248_18, 
        p_wishbone_bd_ram_mem2_248_19, p_wishbone_bd_ram_mem2_248_20, 
        p_wishbone_bd_ram_mem2_248_21, p_wishbone_bd_ram_mem2_248_22, 
        p_wishbone_bd_ram_mem2_248_23, p_wishbone_bd_ram_mem2_249_16, 
        p_wishbone_bd_ram_mem2_249_17, p_wishbone_bd_ram_mem2_249_18, 
        p_wishbone_bd_ram_mem2_249_19, p_wishbone_bd_ram_mem2_249_20, 
        p_wishbone_bd_ram_mem2_249_21, p_wishbone_bd_ram_mem2_249_22, 
        p_wishbone_bd_ram_mem2_249_23, p_wishbone_bd_ram_mem2_250_16, 
        p_wishbone_bd_ram_mem2_250_17, p_wishbone_bd_ram_mem2_250_18, 
        p_wishbone_bd_ram_mem2_250_19, p_wishbone_bd_ram_mem2_250_20, 
        p_wishbone_bd_ram_mem2_250_21, p_wishbone_bd_ram_mem2_250_22, 
        p_wishbone_bd_ram_mem2_250_23, p_wishbone_bd_ram_mem2_251_16, 
        p_wishbone_bd_ram_mem2_251_17, p_wishbone_bd_ram_mem2_251_18, 
        p_wishbone_bd_ram_mem2_251_19, p_wishbone_bd_ram_mem2_251_20, 
        p_wishbone_bd_ram_mem2_251_21, p_wishbone_bd_ram_mem2_251_22, 
        p_wishbone_bd_ram_mem2_251_23, p_wishbone_bd_ram_mem2_252_16, 
        p_wishbone_bd_ram_mem2_252_17, p_wishbone_bd_ram_mem2_252_18, 
        p_wishbone_bd_ram_mem2_252_19, p_wishbone_bd_ram_mem2_252_20, 
        p_wishbone_bd_ram_mem2_252_21, p_wishbone_bd_ram_mem2_252_22, 
        p_wishbone_bd_ram_mem2_252_23, p_wishbone_bd_ram_mem2_253_16, 
        p_wishbone_bd_ram_mem2_253_17, p_wishbone_bd_ram_mem2_253_18, 
        p_wishbone_bd_ram_mem2_253_19, p_wishbone_bd_ram_mem2_253_20, 
        p_wishbone_bd_ram_mem2_253_21, p_wishbone_bd_ram_mem2_253_22, 
        p_wishbone_bd_ram_mem2_253_23, p_wishbone_bd_ram_mem2_254_16, 
        p_wishbone_bd_ram_mem2_254_17, p_wishbone_bd_ram_mem2_254_18, 
        p_wishbone_bd_ram_mem2_254_19, p_wishbone_bd_ram_mem2_254_20, 
        p_wishbone_bd_ram_mem2_254_21, p_wishbone_bd_ram_mem2_254_22, 
        p_wishbone_bd_ram_mem2_254_23, p_wishbone_bd_ram_mem2_255_16, 
        p_wishbone_bd_ram_mem2_255_17, p_wishbone_bd_ram_mem2_255_18, 
        p_wishbone_bd_ram_mem2_255_19, p_wishbone_bd_ram_mem2_255_20, 
        p_wishbone_bd_ram_mem2_255_21, p_wishbone_bd_ram_mem2_255_22, 
        p_wishbone_bd_ram_mem2_255_23, p_wishbone_bd_ram_mem3_0_24, 
        p_wishbone_bd_ram_mem3_0_25, p_wishbone_bd_ram_mem3_0_26, 
        p_wishbone_bd_ram_mem3_0_27, p_wishbone_bd_ram_mem3_0_28, 
        p_wishbone_bd_ram_mem3_0_29, p_wishbone_bd_ram_mem3_0_30, 
        p_wishbone_bd_ram_mem3_0_31, p_wishbone_bd_ram_mem3_1_24, 
        p_wishbone_bd_ram_mem3_1_25, p_wishbone_bd_ram_mem3_1_26, 
        p_wishbone_bd_ram_mem3_1_27, p_wishbone_bd_ram_mem3_1_28, 
        p_wishbone_bd_ram_mem3_1_29, p_wishbone_bd_ram_mem3_1_30, 
        p_wishbone_bd_ram_mem3_1_31, p_wishbone_bd_ram_mem3_2_24, 
        p_wishbone_bd_ram_mem3_2_25, p_wishbone_bd_ram_mem3_2_26, 
        p_wishbone_bd_ram_mem3_2_27, p_wishbone_bd_ram_mem3_2_28, 
        p_wishbone_bd_ram_mem3_2_29, p_wishbone_bd_ram_mem3_2_30, 
        p_wishbone_bd_ram_mem3_2_31, p_wishbone_bd_ram_mem3_3_24, 
        p_wishbone_bd_ram_mem3_3_25, p_wishbone_bd_ram_mem3_3_26, 
        p_wishbone_bd_ram_mem3_3_27, p_wishbone_bd_ram_mem3_3_28, 
        p_wishbone_bd_ram_mem3_3_29, p_wishbone_bd_ram_mem3_3_30, 
        p_wishbone_bd_ram_mem3_3_31, p_wishbone_bd_ram_mem3_4_24, 
        p_wishbone_bd_ram_mem3_4_25, p_wishbone_bd_ram_mem3_4_26, 
        p_wishbone_bd_ram_mem3_4_27, p_wishbone_bd_ram_mem3_4_28, 
        p_wishbone_bd_ram_mem3_4_29, p_wishbone_bd_ram_mem3_4_30, 
        p_wishbone_bd_ram_mem3_4_31, p_wishbone_bd_ram_mem3_5_24, 
        p_wishbone_bd_ram_mem3_5_25, p_wishbone_bd_ram_mem3_5_26, 
        p_wishbone_bd_ram_mem3_5_27, p_wishbone_bd_ram_mem3_5_28, 
        p_wishbone_bd_ram_mem3_5_29, p_wishbone_bd_ram_mem3_5_30, 
        p_wishbone_bd_ram_mem3_5_31, p_wishbone_bd_ram_mem3_6_24, 
        p_wishbone_bd_ram_mem3_6_25, p_wishbone_bd_ram_mem3_6_26, 
        p_wishbone_bd_ram_mem3_6_27, p_wishbone_bd_ram_mem3_6_28, 
        p_wishbone_bd_ram_mem3_6_29, p_wishbone_bd_ram_mem3_6_30, 
        p_wishbone_bd_ram_mem3_6_31, p_wishbone_bd_ram_mem3_7_24, 
        p_wishbone_bd_ram_mem3_7_25, p_wishbone_bd_ram_mem3_7_26, 
        p_wishbone_bd_ram_mem3_7_27, p_wishbone_bd_ram_mem3_7_28, 
        p_wishbone_bd_ram_mem3_7_29, p_wishbone_bd_ram_mem3_7_30, 
        p_wishbone_bd_ram_mem3_7_31, p_wishbone_bd_ram_mem3_8_24, 
        p_wishbone_bd_ram_mem3_8_25, p_wishbone_bd_ram_mem3_8_26, 
        p_wishbone_bd_ram_mem3_8_27, p_wishbone_bd_ram_mem3_8_28, 
        p_wishbone_bd_ram_mem3_8_29, p_wishbone_bd_ram_mem3_8_30, 
        p_wishbone_bd_ram_mem3_8_31, p_wishbone_bd_ram_mem3_9_24, 
        p_wishbone_bd_ram_mem3_9_25, p_wishbone_bd_ram_mem3_9_26, 
        p_wishbone_bd_ram_mem3_9_27, p_wishbone_bd_ram_mem3_9_28, 
        p_wishbone_bd_ram_mem3_9_29, p_wishbone_bd_ram_mem3_9_30, 
        p_wishbone_bd_ram_mem3_9_31, p_wishbone_bd_ram_mem3_10_24, 
        p_wishbone_bd_ram_mem3_10_25, p_wishbone_bd_ram_mem3_10_26, 
        p_wishbone_bd_ram_mem3_10_27, p_wishbone_bd_ram_mem3_10_28, 
        p_wishbone_bd_ram_mem3_10_29, p_wishbone_bd_ram_mem3_10_30, 
        p_wishbone_bd_ram_mem3_10_31, p_wishbone_bd_ram_mem3_11_24, 
        p_wishbone_bd_ram_mem3_11_25, p_wishbone_bd_ram_mem3_11_26, 
        p_wishbone_bd_ram_mem3_11_27, p_wishbone_bd_ram_mem3_11_28, 
        p_wishbone_bd_ram_mem3_11_29, p_wishbone_bd_ram_mem3_11_30, 
        p_wishbone_bd_ram_mem3_11_31, p_wishbone_bd_ram_mem3_12_24, 
        p_wishbone_bd_ram_mem3_12_25, p_wishbone_bd_ram_mem3_12_26, 
        p_wishbone_bd_ram_mem3_12_27, p_wishbone_bd_ram_mem3_12_28, 
        p_wishbone_bd_ram_mem3_12_29, p_wishbone_bd_ram_mem3_12_30, 
        p_wishbone_bd_ram_mem3_12_31, p_wishbone_bd_ram_mem3_13_24, 
        p_wishbone_bd_ram_mem3_13_25, p_wishbone_bd_ram_mem3_13_26, 
        p_wishbone_bd_ram_mem3_13_27, p_wishbone_bd_ram_mem3_13_28, 
        p_wishbone_bd_ram_mem3_13_29, p_wishbone_bd_ram_mem3_13_30, 
        p_wishbone_bd_ram_mem3_13_31, p_wishbone_bd_ram_mem3_14_24, 
        p_wishbone_bd_ram_mem3_14_25, p_wishbone_bd_ram_mem3_14_26, 
        p_wishbone_bd_ram_mem3_14_27, p_wishbone_bd_ram_mem3_14_28, 
        p_wishbone_bd_ram_mem3_14_29, p_wishbone_bd_ram_mem3_14_30, 
        p_wishbone_bd_ram_mem3_14_31, p_wishbone_bd_ram_mem3_15_24, 
        p_wishbone_bd_ram_mem3_15_25, p_wishbone_bd_ram_mem3_15_26, 
        p_wishbone_bd_ram_mem3_15_27, p_wishbone_bd_ram_mem3_15_28, 
        p_wishbone_bd_ram_mem3_15_29, p_wishbone_bd_ram_mem3_15_30, 
        p_wishbone_bd_ram_mem3_15_31, p_wishbone_bd_ram_mem3_16_24, 
        p_wishbone_bd_ram_mem3_16_25, p_wishbone_bd_ram_mem3_16_26, 
        p_wishbone_bd_ram_mem3_16_27, p_wishbone_bd_ram_mem3_16_28, 
        p_wishbone_bd_ram_mem3_16_29, p_wishbone_bd_ram_mem3_16_30, 
        p_wishbone_bd_ram_mem3_16_31, p_wishbone_bd_ram_mem3_17_24, 
        p_wishbone_bd_ram_mem3_17_25, p_wishbone_bd_ram_mem3_17_26, 
        p_wishbone_bd_ram_mem3_17_27, p_wishbone_bd_ram_mem3_17_28, 
        p_wishbone_bd_ram_mem3_17_29, p_wishbone_bd_ram_mem3_17_30, 
        p_wishbone_bd_ram_mem3_17_31, p_wishbone_bd_ram_mem3_18_24, 
        p_wishbone_bd_ram_mem3_18_25, p_wishbone_bd_ram_mem3_18_26, 
        p_wishbone_bd_ram_mem3_18_27, p_wishbone_bd_ram_mem3_18_28, 
        p_wishbone_bd_ram_mem3_18_29, p_wishbone_bd_ram_mem3_18_30, 
        p_wishbone_bd_ram_mem3_18_31, p_wishbone_bd_ram_mem3_19_24, 
        p_wishbone_bd_ram_mem3_19_25, p_wishbone_bd_ram_mem3_19_26, 
        p_wishbone_bd_ram_mem3_19_27, p_wishbone_bd_ram_mem3_19_28, 
        p_wishbone_bd_ram_mem3_19_29, p_wishbone_bd_ram_mem3_19_30, 
        p_wishbone_bd_ram_mem3_19_31, p_wishbone_bd_ram_mem3_20_24, 
        p_wishbone_bd_ram_mem3_20_25, p_wishbone_bd_ram_mem3_20_26, 
        p_wishbone_bd_ram_mem3_20_27, p_wishbone_bd_ram_mem3_20_28, 
        p_wishbone_bd_ram_mem3_20_29, p_wishbone_bd_ram_mem3_20_30, 
        p_wishbone_bd_ram_mem3_20_31, p_wishbone_bd_ram_mem3_21_24, 
        p_wishbone_bd_ram_mem3_21_25, p_wishbone_bd_ram_mem3_21_26, 
        p_wishbone_bd_ram_mem3_21_27, p_wishbone_bd_ram_mem3_21_28, 
        p_wishbone_bd_ram_mem3_21_29, p_wishbone_bd_ram_mem3_21_30, 
        p_wishbone_bd_ram_mem3_21_31, p_wishbone_bd_ram_mem3_22_24, 
        p_wishbone_bd_ram_mem3_22_25, p_wishbone_bd_ram_mem3_22_26, 
        p_wishbone_bd_ram_mem3_22_27, p_wishbone_bd_ram_mem3_22_28, 
        p_wishbone_bd_ram_mem3_22_29, p_wishbone_bd_ram_mem3_22_30, 
        p_wishbone_bd_ram_mem3_22_31, p_wishbone_bd_ram_mem3_23_24, 
        p_wishbone_bd_ram_mem3_23_25, p_wishbone_bd_ram_mem3_23_26, 
        p_wishbone_bd_ram_mem3_23_27, p_wishbone_bd_ram_mem3_23_28, 
        p_wishbone_bd_ram_mem3_23_29, p_wishbone_bd_ram_mem3_23_30, 
        p_wishbone_bd_ram_mem3_23_31, p_wishbone_bd_ram_mem3_24_24, 
        p_wishbone_bd_ram_mem3_24_25, p_wishbone_bd_ram_mem3_24_26, 
        p_wishbone_bd_ram_mem3_24_27, p_wishbone_bd_ram_mem3_24_28, 
        p_wishbone_bd_ram_mem3_24_29, p_wishbone_bd_ram_mem3_24_30, 
        p_wishbone_bd_ram_mem3_24_31, p_wishbone_bd_ram_mem3_25_24, 
        p_wishbone_bd_ram_mem3_25_25, p_wishbone_bd_ram_mem3_25_26, 
        p_wishbone_bd_ram_mem3_25_27, p_wishbone_bd_ram_mem3_25_28, 
        p_wishbone_bd_ram_mem3_25_29, p_wishbone_bd_ram_mem3_25_30, 
        p_wishbone_bd_ram_mem3_25_31, p_wishbone_bd_ram_mem3_26_24, 
        p_wishbone_bd_ram_mem3_26_25, p_wishbone_bd_ram_mem3_26_26, 
        p_wishbone_bd_ram_mem3_26_27, p_wishbone_bd_ram_mem3_26_28, 
        p_wishbone_bd_ram_mem3_26_29, p_wishbone_bd_ram_mem3_26_30, 
        p_wishbone_bd_ram_mem3_26_31, p_wishbone_bd_ram_mem3_27_24, 
        p_wishbone_bd_ram_mem3_27_25, p_wishbone_bd_ram_mem3_27_26, 
        p_wishbone_bd_ram_mem3_27_27, p_wishbone_bd_ram_mem3_27_28, 
        p_wishbone_bd_ram_mem3_27_29, p_wishbone_bd_ram_mem3_27_30, 
        p_wishbone_bd_ram_mem3_27_31, p_wishbone_bd_ram_mem3_28_24, 
        p_wishbone_bd_ram_mem3_28_25, p_wishbone_bd_ram_mem3_28_26, 
        p_wishbone_bd_ram_mem3_28_27, p_wishbone_bd_ram_mem3_28_28, 
        p_wishbone_bd_ram_mem3_28_29, p_wishbone_bd_ram_mem3_28_30, 
        p_wishbone_bd_ram_mem3_28_31, p_wishbone_bd_ram_mem3_29_24, 
        p_wishbone_bd_ram_mem3_29_25, p_wishbone_bd_ram_mem3_29_26, 
        p_wishbone_bd_ram_mem3_29_27, p_wishbone_bd_ram_mem3_29_28, 
        p_wishbone_bd_ram_mem3_29_29, p_wishbone_bd_ram_mem3_29_30, 
        p_wishbone_bd_ram_mem3_29_31, p_wishbone_bd_ram_mem3_30_24, 
        p_wishbone_bd_ram_mem3_30_25, p_wishbone_bd_ram_mem3_30_26, 
        p_wishbone_bd_ram_mem3_30_27, p_wishbone_bd_ram_mem3_30_28, 
        p_wishbone_bd_ram_mem3_30_29, p_wishbone_bd_ram_mem3_30_30, 
        p_wishbone_bd_ram_mem3_30_31, p_wishbone_bd_ram_mem3_31_24, 
        p_wishbone_bd_ram_mem3_31_25, p_wishbone_bd_ram_mem3_31_26, 
        p_wishbone_bd_ram_mem3_31_27, p_wishbone_bd_ram_mem3_31_28, 
        p_wishbone_bd_ram_mem3_31_29, p_wishbone_bd_ram_mem3_31_30, 
        p_wishbone_bd_ram_mem3_31_31, p_wishbone_bd_ram_mem3_32_24, 
        p_wishbone_bd_ram_mem3_32_25, p_wishbone_bd_ram_mem3_32_26, 
        p_wishbone_bd_ram_mem3_32_27, p_wishbone_bd_ram_mem3_32_28, 
        p_wishbone_bd_ram_mem3_32_29, p_wishbone_bd_ram_mem3_32_30, 
        p_wishbone_bd_ram_mem3_32_31, p_wishbone_bd_ram_mem3_33_24, 
        p_wishbone_bd_ram_mem3_33_25, p_wishbone_bd_ram_mem3_33_26, 
        p_wishbone_bd_ram_mem3_33_27, p_wishbone_bd_ram_mem3_33_28, 
        p_wishbone_bd_ram_mem3_33_29, p_wishbone_bd_ram_mem3_33_30, 
        p_wishbone_bd_ram_mem3_33_31, p_wishbone_bd_ram_mem3_34_24, 
        p_wishbone_bd_ram_mem3_34_25, p_wishbone_bd_ram_mem3_34_26, 
        p_wishbone_bd_ram_mem3_34_27, p_wishbone_bd_ram_mem3_34_28, 
        p_wishbone_bd_ram_mem3_34_29, p_wishbone_bd_ram_mem3_34_30, 
        p_wishbone_bd_ram_mem3_34_31, p_wishbone_bd_ram_mem3_35_24, 
        p_wishbone_bd_ram_mem3_35_25, p_wishbone_bd_ram_mem3_35_26, 
        p_wishbone_bd_ram_mem3_35_27, p_wishbone_bd_ram_mem3_35_28, 
        p_wishbone_bd_ram_mem3_35_29, p_wishbone_bd_ram_mem3_35_30, 
        p_wishbone_bd_ram_mem3_35_31, p_wishbone_bd_ram_mem3_36_24, 
        p_wishbone_bd_ram_mem3_36_25, p_wishbone_bd_ram_mem3_36_26, 
        p_wishbone_bd_ram_mem3_36_27, p_wishbone_bd_ram_mem3_36_28, 
        p_wishbone_bd_ram_mem3_36_29, p_wishbone_bd_ram_mem3_36_30, 
        p_wishbone_bd_ram_mem3_36_31, p_wishbone_bd_ram_mem3_37_24, 
        p_wishbone_bd_ram_mem3_37_25, p_wishbone_bd_ram_mem3_37_26, 
        p_wishbone_bd_ram_mem3_37_27, p_wishbone_bd_ram_mem3_37_28, 
        p_wishbone_bd_ram_mem3_37_29, p_wishbone_bd_ram_mem3_37_30, 
        p_wishbone_bd_ram_mem3_37_31, p_wishbone_bd_ram_mem3_38_24, 
        p_wishbone_bd_ram_mem3_38_25, p_wishbone_bd_ram_mem3_38_26, 
        p_wishbone_bd_ram_mem3_38_27, p_wishbone_bd_ram_mem3_38_28, 
        p_wishbone_bd_ram_mem3_38_29, p_wishbone_bd_ram_mem3_38_30, 
        p_wishbone_bd_ram_mem3_38_31, p_wishbone_bd_ram_mem3_39_24, 
        p_wishbone_bd_ram_mem3_39_25, p_wishbone_bd_ram_mem3_39_26, 
        p_wishbone_bd_ram_mem3_39_27, p_wishbone_bd_ram_mem3_39_28, 
        p_wishbone_bd_ram_mem3_39_29, p_wishbone_bd_ram_mem3_39_30, 
        p_wishbone_bd_ram_mem3_39_31, p_wishbone_bd_ram_mem3_40_24, 
        p_wishbone_bd_ram_mem3_40_25, p_wishbone_bd_ram_mem3_40_26, 
        p_wishbone_bd_ram_mem3_40_27, p_wishbone_bd_ram_mem3_40_28, 
        p_wishbone_bd_ram_mem3_40_29, p_wishbone_bd_ram_mem3_40_30, 
        p_wishbone_bd_ram_mem3_40_31, p_wishbone_bd_ram_mem3_41_24, 
        p_wishbone_bd_ram_mem3_41_25, p_wishbone_bd_ram_mem3_41_26, 
        p_wishbone_bd_ram_mem3_41_27, p_wishbone_bd_ram_mem3_41_28, 
        p_wishbone_bd_ram_mem3_41_29, p_wishbone_bd_ram_mem3_41_30, 
        p_wishbone_bd_ram_mem3_41_31, p_wishbone_bd_ram_mem3_42_24, 
        p_wishbone_bd_ram_mem3_42_25, p_wishbone_bd_ram_mem3_42_26, 
        p_wishbone_bd_ram_mem3_42_27, p_wishbone_bd_ram_mem3_42_28, 
        p_wishbone_bd_ram_mem3_42_29, p_wishbone_bd_ram_mem3_42_30, 
        p_wishbone_bd_ram_mem3_42_31, p_wishbone_bd_ram_mem3_43_24, 
        p_wishbone_bd_ram_mem3_43_25, p_wishbone_bd_ram_mem3_43_26, 
        p_wishbone_bd_ram_mem3_43_27, p_wishbone_bd_ram_mem3_43_28, 
        p_wishbone_bd_ram_mem3_43_29, p_wishbone_bd_ram_mem3_43_30, 
        p_wishbone_bd_ram_mem3_43_31, p_wishbone_bd_ram_mem3_44_24, 
        p_wishbone_bd_ram_mem3_44_25, p_wishbone_bd_ram_mem3_44_26, 
        p_wishbone_bd_ram_mem3_44_27, p_wishbone_bd_ram_mem3_44_28, 
        p_wishbone_bd_ram_mem3_44_29, p_wishbone_bd_ram_mem3_44_30, 
        p_wishbone_bd_ram_mem3_44_31, p_wishbone_bd_ram_mem3_45_24, 
        p_wishbone_bd_ram_mem3_45_25, p_wishbone_bd_ram_mem3_45_26, 
        p_wishbone_bd_ram_mem3_45_27, p_wishbone_bd_ram_mem3_45_28, 
        p_wishbone_bd_ram_mem3_45_29, p_wishbone_bd_ram_mem3_45_30, 
        p_wishbone_bd_ram_mem3_45_31, p_wishbone_bd_ram_mem3_46_24, 
        p_wishbone_bd_ram_mem3_46_25, p_wishbone_bd_ram_mem3_46_26, 
        p_wishbone_bd_ram_mem3_46_27, p_wishbone_bd_ram_mem3_46_28, 
        p_wishbone_bd_ram_mem3_46_29, p_wishbone_bd_ram_mem3_46_30, 
        p_wishbone_bd_ram_mem3_46_31, p_wishbone_bd_ram_mem3_47_24, 
        p_wishbone_bd_ram_mem3_47_25, p_wishbone_bd_ram_mem3_47_26, 
        p_wishbone_bd_ram_mem3_47_27, p_wishbone_bd_ram_mem3_47_28, 
        p_wishbone_bd_ram_mem3_47_29, p_wishbone_bd_ram_mem3_47_30, 
        p_wishbone_bd_ram_mem3_47_31, p_wishbone_bd_ram_mem3_48_24, 
        p_wishbone_bd_ram_mem3_48_25, p_wishbone_bd_ram_mem3_48_26, 
        p_wishbone_bd_ram_mem3_48_27, p_wishbone_bd_ram_mem3_48_28, 
        p_wishbone_bd_ram_mem3_48_29, p_wishbone_bd_ram_mem3_48_30, 
        p_wishbone_bd_ram_mem3_48_31, p_wishbone_bd_ram_mem3_49_24, 
        p_wishbone_bd_ram_mem3_49_25, p_wishbone_bd_ram_mem3_49_26, 
        p_wishbone_bd_ram_mem3_49_27, p_wishbone_bd_ram_mem3_49_28, 
        p_wishbone_bd_ram_mem3_49_29, p_wishbone_bd_ram_mem3_49_30, 
        p_wishbone_bd_ram_mem3_49_31, p_wishbone_bd_ram_mem3_50_24, 
        p_wishbone_bd_ram_mem3_50_25, p_wishbone_bd_ram_mem3_50_26, 
        p_wishbone_bd_ram_mem3_50_27, p_wishbone_bd_ram_mem3_50_28, 
        p_wishbone_bd_ram_mem3_50_29, p_wishbone_bd_ram_mem3_50_30, 
        p_wishbone_bd_ram_mem3_50_31, p_wishbone_bd_ram_mem3_51_24, 
        p_wishbone_bd_ram_mem3_51_25, p_wishbone_bd_ram_mem3_51_26, 
        p_wishbone_bd_ram_mem3_51_27, p_wishbone_bd_ram_mem3_51_28, 
        p_wishbone_bd_ram_mem3_51_29, p_wishbone_bd_ram_mem3_51_30, 
        p_wishbone_bd_ram_mem3_51_31, p_wishbone_bd_ram_mem3_52_24, 
        p_wishbone_bd_ram_mem3_52_25, p_wishbone_bd_ram_mem3_52_26, 
        p_wishbone_bd_ram_mem3_52_27, p_wishbone_bd_ram_mem3_52_28, 
        p_wishbone_bd_ram_mem3_52_29, p_wishbone_bd_ram_mem3_52_30, 
        p_wishbone_bd_ram_mem3_52_31, p_wishbone_bd_ram_mem3_53_24, 
        p_wishbone_bd_ram_mem3_53_25, p_wishbone_bd_ram_mem3_53_26, 
        p_wishbone_bd_ram_mem3_53_27, p_wishbone_bd_ram_mem3_53_28, 
        p_wishbone_bd_ram_mem3_53_29, p_wishbone_bd_ram_mem3_53_30, 
        p_wishbone_bd_ram_mem3_53_31, p_wishbone_bd_ram_mem3_54_24, 
        p_wishbone_bd_ram_mem3_54_25, p_wishbone_bd_ram_mem3_54_26, 
        p_wishbone_bd_ram_mem3_54_27, p_wishbone_bd_ram_mem3_54_28, 
        p_wishbone_bd_ram_mem3_54_29, p_wishbone_bd_ram_mem3_54_30, 
        p_wishbone_bd_ram_mem3_54_31, p_wishbone_bd_ram_mem3_55_24, 
        p_wishbone_bd_ram_mem3_55_25, p_wishbone_bd_ram_mem3_55_26, 
        p_wishbone_bd_ram_mem3_55_27, p_wishbone_bd_ram_mem3_55_28, 
        p_wishbone_bd_ram_mem3_55_29, p_wishbone_bd_ram_mem3_55_30, 
        p_wishbone_bd_ram_mem3_55_31, p_wishbone_bd_ram_mem3_56_24, 
        p_wishbone_bd_ram_mem3_56_25, p_wishbone_bd_ram_mem3_56_26, 
        p_wishbone_bd_ram_mem3_56_27, p_wishbone_bd_ram_mem3_56_28, 
        p_wishbone_bd_ram_mem3_56_29, p_wishbone_bd_ram_mem3_56_30, 
        p_wishbone_bd_ram_mem3_56_31, p_wishbone_bd_ram_mem3_57_24, 
        p_wishbone_bd_ram_mem3_57_25, p_wishbone_bd_ram_mem3_57_26, 
        p_wishbone_bd_ram_mem3_57_27, p_wishbone_bd_ram_mem3_57_28, 
        p_wishbone_bd_ram_mem3_57_29, p_wishbone_bd_ram_mem3_57_30, 
        p_wishbone_bd_ram_mem3_57_31, p_wishbone_bd_ram_mem3_58_24, 
        p_wishbone_bd_ram_mem3_58_25, p_wishbone_bd_ram_mem3_58_26, 
        p_wishbone_bd_ram_mem3_58_27, p_wishbone_bd_ram_mem3_58_28, 
        p_wishbone_bd_ram_mem3_58_29, p_wishbone_bd_ram_mem3_58_30, 
        p_wishbone_bd_ram_mem3_58_31, p_wishbone_bd_ram_mem3_59_24, 
        p_wishbone_bd_ram_mem3_59_25, p_wishbone_bd_ram_mem3_59_26, 
        p_wishbone_bd_ram_mem3_59_27, p_wishbone_bd_ram_mem3_59_28, 
        p_wishbone_bd_ram_mem3_59_29, p_wishbone_bd_ram_mem3_59_30, 
        p_wishbone_bd_ram_mem3_59_31, p_wishbone_bd_ram_mem3_60_24, 
        p_wishbone_bd_ram_mem3_60_25, p_wishbone_bd_ram_mem3_60_26, 
        p_wishbone_bd_ram_mem3_60_27, p_wishbone_bd_ram_mem3_60_28, 
        p_wishbone_bd_ram_mem3_60_29, p_wishbone_bd_ram_mem3_60_30, 
        p_wishbone_bd_ram_mem3_60_31, p_wishbone_bd_ram_mem3_61_24, 
        p_wishbone_bd_ram_mem3_61_25, p_wishbone_bd_ram_mem3_61_26, 
        p_wishbone_bd_ram_mem3_61_27, p_wishbone_bd_ram_mem3_61_28, 
        p_wishbone_bd_ram_mem3_61_29, p_wishbone_bd_ram_mem3_61_30, 
        p_wishbone_bd_ram_mem3_61_31, p_wishbone_bd_ram_mem3_62_24, 
        p_wishbone_bd_ram_mem3_62_25, p_wishbone_bd_ram_mem3_62_26, 
        p_wishbone_bd_ram_mem3_62_27, p_wishbone_bd_ram_mem3_62_28, 
        p_wishbone_bd_ram_mem3_62_29, p_wishbone_bd_ram_mem3_62_30, 
        p_wishbone_bd_ram_mem3_62_31, p_wishbone_bd_ram_mem3_63_24, 
        p_wishbone_bd_ram_mem3_63_25, p_wishbone_bd_ram_mem3_63_26, 
        p_wishbone_bd_ram_mem3_63_27, p_wishbone_bd_ram_mem3_63_28, 
        p_wishbone_bd_ram_mem3_63_29, p_wishbone_bd_ram_mem3_63_30, 
        p_wishbone_bd_ram_mem3_63_31, p_wishbone_bd_ram_mem3_64_24, 
        p_wishbone_bd_ram_mem3_64_25, p_wishbone_bd_ram_mem3_64_26, 
        p_wishbone_bd_ram_mem3_64_27, p_wishbone_bd_ram_mem3_64_28, 
        p_wishbone_bd_ram_mem3_64_29, p_wishbone_bd_ram_mem3_64_30, 
        p_wishbone_bd_ram_mem3_64_31, p_wishbone_bd_ram_mem3_65_24, 
        p_wishbone_bd_ram_mem3_65_25, p_wishbone_bd_ram_mem3_65_26, 
        p_wishbone_bd_ram_mem3_65_27, p_wishbone_bd_ram_mem3_65_28, 
        p_wishbone_bd_ram_mem3_65_29, p_wishbone_bd_ram_mem3_65_30, 
        p_wishbone_bd_ram_mem3_65_31, p_wishbone_bd_ram_mem3_66_24, 
        p_wishbone_bd_ram_mem3_66_25, p_wishbone_bd_ram_mem3_66_26, 
        p_wishbone_bd_ram_mem3_66_27, p_wishbone_bd_ram_mem3_66_28, 
        p_wishbone_bd_ram_mem3_66_29, p_wishbone_bd_ram_mem3_66_30, 
        p_wishbone_bd_ram_mem3_66_31, p_wishbone_bd_ram_mem3_67_24, 
        p_wishbone_bd_ram_mem3_67_25, p_wishbone_bd_ram_mem3_67_26, 
        p_wishbone_bd_ram_mem3_67_27, p_wishbone_bd_ram_mem3_67_28, 
        p_wishbone_bd_ram_mem3_67_29, p_wishbone_bd_ram_mem3_67_30, 
        p_wishbone_bd_ram_mem3_67_31, p_wishbone_bd_ram_mem3_68_24, 
        p_wishbone_bd_ram_mem3_68_25, p_wishbone_bd_ram_mem3_68_26, 
        p_wishbone_bd_ram_mem3_68_27, p_wishbone_bd_ram_mem3_68_28, 
        p_wishbone_bd_ram_mem3_68_29, p_wishbone_bd_ram_mem3_68_30, 
        p_wishbone_bd_ram_mem3_68_31, p_wishbone_bd_ram_mem3_69_24, 
        p_wishbone_bd_ram_mem3_69_25, p_wishbone_bd_ram_mem3_69_26, 
        p_wishbone_bd_ram_mem3_69_27, p_wishbone_bd_ram_mem3_69_28, 
        p_wishbone_bd_ram_mem3_69_29, p_wishbone_bd_ram_mem3_69_30, 
        p_wishbone_bd_ram_mem3_69_31, p_wishbone_bd_ram_mem3_70_24, 
        p_wishbone_bd_ram_mem3_70_25, p_wishbone_bd_ram_mem3_70_26, 
        p_wishbone_bd_ram_mem3_70_27, p_wishbone_bd_ram_mem3_70_28, 
        p_wishbone_bd_ram_mem3_70_29, p_wishbone_bd_ram_mem3_70_30, 
        p_wishbone_bd_ram_mem3_70_31, p_wishbone_bd_ram_mem3_71_24, 
        p_wishbone_bd_ram_mem3_71_25, p_wishbone_bd_ram_mem3_71_26, 
        p_wishbone_bd_ram_mem3_71_27, p_wishbone_bd_ram_mem3_71_28, 
        p_wishbone_bd_ram_mem3_71_29, p_wishbone_bd_ram_mem3_71_30, 
        p_wishbone_bd_ram_mem3_71_31, p_wishbone_bd_ram_mem3_72_24, 
        p_wishbone_bd_ram_mem3_72_25, p_wishbone_bd_ram_mem3_72_26, 
        p_wishbone_bd_ram_mem3_72_27, p_wishbone_bd_ram_mem3_72_28, 
        p_wishbone_bd_ram_mem3_72_29, p_wishbone_bd_ram_mem3_72_30, 
        p_wishbone_bd_ram_mem3_72_31, p_wishbone_bd_ram_mem3_73_24, 
        p_wishbone_bd_ram_mem3_73_25, p_wishbone_bd_ram_mem3_73_26, 
        p_wishbone_bd_ram_mem3_73_27, p_wishbone_bd_ram_mem3_73_28, 
        p_wishbone_bd_ram_mem3_73_29, p_wishbone_bd_ram_mem3_73_30, 
        p_wishbone_bd_ram_mem3_73_31, p_wishbone_bd_ram_mem3_74_24, 
        p_wishbone_bd_ram_mem3_74_25, p_wishbone_bd_ram_mem3_74_26, 
        p_wishbone_bd_ram_mem3_74_27, p_wishbone_bd_ram_mem3_74_28, 
        p_wishbone_bd_ram_mem3_74_29, p_wishbone_bd_ram_mem3_74_30, 
        p_wishbone_bd_ram_mem3_74_31, p_wishbone_bd_ram_mem3_75_24, 
        p_wishbone_bd_ram_mem3_75_25, p_wishbone_bd_ram_mem3_75_26, 
        p_wishbone_bd_ram_mem3_75_27, p_wishbone_bd_ram_mem3_75_28, 
        p_wishbone_bd_ram_mem3_75_29, p_wishbone_bd_ram_mem3_75_30, 
        p_wishbone_bd_ram_mem3_75_31, p_wishbone_bd_ram_mem3_76_24, 
        p_wishbone_bd_ram_mem3_76_25, p_wishbone_bd_ram_mem3_76_26, 
        p_wishbone_bd_ram_mem3_76_27, p_wishbone_bd_ram_mem3_76_28, 
        p_wishbone_bd_ram_mem3_76_29, p_wishbone_bd_ram_mem3_76_30, 
        p_wishbone_bd_ram_mem3_76_31, p_wishbone_bd_ram_mem3_77_24, 
        p_wishbone_bd_ram_mem3_77_25, p_wishbone_bd_ram_mem3_77_26, 
        p_wishbone_bd_ram_mem3_77_27, p_wishbone_bd_ram_mem3_77_28, 
        p_wishbone_bd_ram_mem3_77_29, p_wishbone_bd_ram_mem3_77_30, 
        p_wishbone_bd_ram_mem3_77_31, p_wishbone_bd_ram_mem3_78_24, 
        p_wishbone_bd_ram_mem3_78_25, p_wishbone_bd_ram_mem3_78_26, 
        p_wishbone_bd_ram_mem3_78_27, p_wishbone_bd_ram_mem3_78_28, 
        p_wishbone_bd_ram_mem3_78_29, p_wishbone_bd_ram_mem3_78_30, 
        p_wishbone_bd_ram_mem3_78_31, p_wishbone_bd_ram_mem3_79_24, 
        p_wishbone_bd_ram_mem3_79_25, p_wishbone_bd_ram_mem3_79_26, 
        p_wishbone_bd_ram_mem3_79_27, p_wishbone_bd_ram_mem3_79_28, 
        p_wishbone_bd_ram_mem3_79_29, p_wishbone_bd_ram_mem3_79_30, 
        p_wishbone_bd_ram_mem3_79_31, p_wishbone_bd_ram_mem3_80_24, 
        p_wishbone_bd_ram_mem3_80_25, p_wishbone_bd_ram_mem3_80_26, 
        p_wishbone_bd_ram_mem3_80_27, p_wishbone_bd_ram_mem3_80_28, 
        p_wishbone_bd_ram_mem3_80_29, p_wishbone_bd_ram_mem3_80_30, 
        p_wishbone_bd_ram_mem3_80_31, p_wishbone_bd_ram_mem3_81_24, 
        p_wishbone_bd_ram_mem3_81_25, p_wishbone_bd_ram_mem3_81_26, 
        p_wishbone_bd_ram_mem3_81_27, p_wishbone_bd_ram_mem3_81_28, 
        p_wishbone_bd_ram_mem3_81_29, p_wishbone_bd_ram_mem3_81_30, 
        p_wishbone_bd_ram_mem3_81_31, p_wishbone_bd_ram_mem3_82_24, 
        p_wishbone_bd_ram_mem3_82_25, p_wishbone_bd_ram_mem3_82_26, 
        p_wishbone_bd_ram_mem3_82_27, p_wishbone_bd_ram_mem3_82_28, 
        p_wishbone_bd_ram_mem3_82_29, p_wishbone_bd_ram_mem3_82_30, 
        p_wishbone_bd_ram_mem3_82_31, p_wishbone_bd_ram_mem3_83_24, 
        p_wishbone_bd_ram_mem3_83_25, p_wishbone_bd_ram_mem3_83_26, 
        p_wishbone_bd_ram_mem3_83_27, p_wishbone_bd_ram_mem3_83_28, 
        p_wishbone_bd_ram_mem3_83_29, p_wishbone_bd_ram_mem3_83_30, 
        p_wishbone_bd_ram_mem3_83_31, p_wishbone_bd_ram_mem3_84_24, 
        p_wishbone_bd_ram_mem3_84_25, p_wishbone_bd_ram_mem3_84_26, 
        p_wishbone_bd_ram_mem3_84_27, p_wishbone_bd_ram_mem3_84_28, 
        p_wishbone_bd_ram_mem3_84_29, p_wishbone_bd_ram_mem3_84_30, 
        p_wishbone_bd_ram_mem3_84_31, p_wishbone_bd_ram_mem3_85_24, 
        p_wishbone_bd_ram_mem3_85_25, p_wishbone_bd_ram_mem3_85_26, 
        p_wishbone_bd_ram_mem3_85_27, p_wishbone_bd_ram_mem3_85_28, 
        p_wishbone_bd_ram_mem3_85_29, p_wishbone_bd_ram_mem3_85_30, 
        p_wishbone_bd_ram_mem3_85_31, p_wishbone_bd_ram_mem3_86_24, 
        p_wishbone_bd_ram_mem3_86_25, p_wishbone_bd_ram_mem3_86_26, 
        p_wishbone_bd_ram_mem3_86_27, p_wishbone_bd_ram_mem3_86_28, 
        p_wishbone_bd_ram_mem3_86_29, p_wishbone_bd_ram_mem3_86_30, 
        p_wishbone_bd_ram_mem3_86_31, p_wishbone_bd_ram_mem3_87_24, 
        p_wishbone_bd_ram_mem3_87_25, p_wishbone_bd_ram_mem3_87_26, 
        p_wishbone_bd_ram_mem3_87_27, p_wishbone_bd_ram_mem3_87_28, 
        p_wishbone_bd_ram_mem3_87_29, p_wishbone_bd_ram_mem3_87_30, 
        p_wishbone_bd_ram_mem3_87_31, p_wishbone_bd_ram_mem3_88_24, 
        p_wishbone_bd_ram_mem3_88_25, p_wishbone_bd_ram_mem3_88_26, 
        p_wishbone_bd_ram_mem3_88_27, p_wishbone_bd_ram_mem3_88_28, 
        p_wishbone_bd_ram_mem3_88_29, p_wishbone_bd_ram_mem3_88_30, 
        p_wishbone_bd_ram_mem3_88_31, p_wishbone_bd_ram_mem3_89_24, 
        p_wishbone_bd_ram_mem3_89_25, p_wishbone_bd_ram_mem3_89_26, 
        p_wishbone_bd_ram_mem3_89_27, p_wishbone_bd_ram_mem3_89_28, 
        p_wishbone_bd_ram_mem3_89_29, p_wishbone_bd_ram_mem3_89_30, 
        p_wishbone_bd_ram_mem3_89_31, p_wishbone_bd_ram_mem3_90_24, 
        p_wishbone_bd_ram_mem3_90_25, p_wishbone_bd_ram_mem3_90_26, 
        p_wishbone_bd_ram_mem3_90_27, p_wishbone_bd_ram_mem3_90_28, 
        p_wishbone_bd_ram_mem3_90_29, p_wishbone_bd_ram_mem3_90_30, 
        p_wishbone_bd_ram_mem3_90_31, p_wishbone_bd_ram_mem3_91_24, 
        p_wishbone_bd_ram_mem3_91_25, p_wishbone_bd_ram_mem3_91_26, 
        p_wishbone_bd_ram_mem3_91_27, p_wishbone_bd_ram_mem3_91_28, 
        p_wishbone_bd_ram_mem3_91_29, p_wishbone_bd_ram_mem3_91_30, 
        p_wishbone_bd_ram_mem3_91_31, p_wishbone_bd_ram_mem3_92_24, 
        p_wishbone_bd_ram_mem3_92_25, p_wishbone_bd_ram_mem3_92_26, 
        p_wishbone_bd_ram_mem3_92_27, p_wishbone_bd_ram_mem3_92_28, 
        p_wishbone_bd_ram_mem3_92_29, p_wishbone_bd_ram_mem3_92_30, 
        p_wishbone_bd_ram_mem3_92_31, p_wishbone_bd_ram_mem3_93_24, 
        p_wishbone_bd_ram_mem3_93_25, p_wishbone_bd_ram_mem3_93_26, 
        p_wishbone_bd_ram_mem3_93_27, p_wishbone_bd_ram_mem3_93_28, 
        p_wishbone_bd_ram_mem3_93_29, p_wishbone_bd_ram_mem3_93_30, 
        p_wishbone_bd_ram_mem3_93_31, p_wishbone_bd_ram_mem3_94_24, 
        p_wishbone_bd_ram_mem3_94_25, p_wishbone_bd_ram_mem3_94_26, 
        p_wishbone_bd_ram_mem3_94_27, p_wishbone_bd_ram_mem3_94_28, 
        p_wishbone_bd_ram_mem3_94_29, p_wishbone_bd_ram_mem3_94_30, 
        p_wishbone_bd_ram_mem3_94_31, p_wishbone_bd_ram_mem3_95_24, 
        p_wishbone_bd_ram_mem3_95_25, p_wishbone_bd_ram_mem3_95_26, 
        p_wishbone_bd_ram_mem3_95_27, p_wishbone_bd_ram_mem3_95_28, 
        p_wishbone_bd_ram_mem3_95_29, p_wishbone_bd_ram_mem3_95_30, 
        p_wishbone_bd_ram_mem3_95_31, p_wishbone_bd_ram_mem3_96_24, 
        p_wishbone_bd_ram_mem3_96_25, p_wishbone_bd_ram_mem3_96_26, 
        p_wishbone_bd_ram_mem3_96_27, p_wishbone_bd_ram_mem3_96_28, 
        p_wishbone_bd_ram_mem3_96_29, p_wishbone_bd_ram_mem3_96_30, 
        p_wishbone_bd_ram_mem3_96_31, p_wishbone_bd_ram_mem3_97_24, 
        p_wishbone_bd_ram_mem3_97_25, p_wishbone_bd_ram_mem3_97_26, 
        p_wishbone_bd_ram_mem3_97_27, p_wishbone_bd_ram_mem3_97_28, 
        p_wishbone_bd_ram_mem3_97_29, p_wishbone_bd_ram_mem3_97_30, 
        p_wishbone_bd_ram_mem3_97_31, p_wishbone_bd_ram_mem3_98_24, 
        p_wishbone_bd_ram_mem3_98_25, p_wishbone_bd_ram_mem3_98_26, 
        p_wishbone_bd_ram_mem3_98_27, p_wishbone_bd_ram_mem3_98_28, 
        p_wishbone_bd_ram_mem3_98_29, p_wishbone_bd_ram_mem3_98_30, 
        p_wishbone_bd_ram_mem3_98_31, p_wishbone_bd_ram_mem3_99_24, 
        p_wishbone_bd_ram_mem3_99_25, p_wishbone_bd_ram_mem3_99_26, 
        p_wishbone_bd_ram_mem3_99_27, p_wishbone_bd_ram_mem3_99_28, 
        p_wishbone_bd_ram_mem3_99_29, p_wishbone_bd_ram_mem3_99_30, 
        p_wishbone_bd_ram_mem3_99_31, p_wishbone_bd_ram_mem3_100_24, 
        p_wishbone_bd_ram_mem3_100_25, p_wishbone_bd_ram_mem3_100_26, 
        p_wishbone_bd_ram_mem3_100_27, p_wishbone_bd_ram_mem3_100_28, 
        p_wishbone_bd_ram_mem3_100_29, p_wishbone_bd_ram_mem3_100_30, 
        p_wishbone_bd_ram_mem3_100_31, p_wishbone_bd_ram_mem3_101_24, 
        p_wishbone_bd_ram_mem3_101_25, p_wishbone_bd_ram_mem3_101_26, 
        p_wishbone_bd_ram_mem3_101_27, p_wishbone_bd_ram_mem3_101_28, 
        p_wishbone_bd_ram_mem3_101_29, p_wishbone_bd_ram_mem3_101_30, 
        p_wishbone_bd_ram_mem3_101_31, p_wishbone_bd_ram_mem3_102_24, 
        p_wishbone_bd_ram_mem3_102_25, p_wishbone_bd_ram_mem3_102_26, 
        p_wishbone_bd_ram_mem3_102_27, p_wishbone_bd_ram_mem3_102_28, 
        p_wishbone_bd_ram_mem3_102_29, p_wishbone_bd_ram_mem3_102_30, 
        p_wishbone_bd_ram_mem3_102_31, p_wishbone_bd_ram_mem3_103_24, 
        p_wishbone_bd_ram_mem3_103_25, p_wishbone_bd_ram_mem3_103_26, 
        p_wishbone_bd_ram_mem3_103_27, p_wishbone_bd_ram_mem3_103_28, 
        p_wishbone_bd_ram_mem3_103_29, p_wishbone_bd_ram_mem3_103_30, 
        p_wishbone_bd_ram_mem3_103_31, p_wishbone_bd_ram_mem3_104_24, 
        p_wishbone_bd_ram_mem3_104_25, p_wishbone_bd_ram_mem3_104_26, 
        p_wishbone_bd_ram_mem3_104_27, p_wishbone_bd_ram_mem3_104_28, 
        p_wishbone_bd_ram_mem3_104_29, p_wishbone_bd_ram_mem3_104_30, 
        p_wishbone_bd_ram_mem3_104_31, p_wishbone_bd_ram_mem3_105_24, 
        p_wishbone_bd_ram_mem3_105_25, p_wishbone_bd_ram_mem3_105_26, 
        p_wishbone_bd_ram_mem3_105_27, p_wishbone_bd_ram_mem3_105_28, 
        p_wishbone_bd_ram_mem3_105_29, p_wishbone_bd_ram_mem3_105_30, 
        p_wishbone_bd_ram_mem3_105_31, p_wishbone_bd_ram_mem3_106_24, 
        p_wishbone_bd_ram_mem3_106_25, p_wishbone_bd_ram_mem3_106_26, 
        p_wishbone_bd_ram_mem3_106_27, p_wishbone_bd_ram_mem3_106_28, 
        p_wishbone_bd_ram_mem3_106_29, p_wishbone_bd_ram_mem3_106_30, 
        p_wishbone_bd_ram_mem3_106_31, p_wishbone_bd_ram_mem3_107_24, 
        p_wishbone_bd_ram_mem3_107_25, p_wishbone_bd_ram_mem3_107_26, 
        p_wishbone_bd_ram_mem3_107_27, p_wishbone_bd_ram_mem3_107_28, 
        p_wishbone_bd_ram_mem3_107_29, p_wishbone_bd_ram_mem3_107_30, 
        p_wishbone_bd_ram_mem3_107_31, p_wishbone_bd_ram_mem3_108_24, 
        p_wishbone_bd_ram_mem3_108_25, p_wishbone_bd_ram_mem3_108_26, 
        p_wishbone_bd_ram_mem3_108_27, p_wishbone_bd_ram_mem3_108_28, 
        p_wishbone_bd_ram_mem3_108_29, p_wishbone_bd_ram_mem3_108_30, 
        p_wishbone_bd_ram_mem3_108_31, p_wishbone_bd_ram_mem3_109_24, 
        p_wishbone_bd_ram_mem3_109_25, p_wishbone_bd_ram_mem3_109_26, 
        p_wishbone_bd_ram_mem3_109_27, p_wishbone_bd_ram_mem3_109_28, 
        p_wishbone_bd_ram_mem3_109_29, p_wishbone_bd_ram_mem3_109_30, 
        p_wishbone_bd_ram_mem3_109_31, p_wishbone_bd_ram_mem3_110_24, 
        p_wishbone_bd_ram_mem3_110_25, p_wishbone_bd_ram_mem3_110_26, 
        p_wishbone_bd_ram_mem3_110_27, p_wishbone_bd_ram_mem3_110_28, 
        p_wishbone_bd_ram_mem3_110_29, p_wishbone_bd_ram_mem3_110_30, 
        p_wishbone_bd_ram_mem3_110_31, p_wishbone_bd_ram_mem3_111_24, 
        p_wishbone_bd_ram_mem3_111_25, p_wishbone_bd_ram_mem3_111_26, 
        p_wishbone_bd_ram_mem3_111_27, p_wishbone_bd_ram_mem3_111_28, 
        p_wishbone_bd_ram_mem3_111_29, p_wishbone_bd_ram_mem3_111_30, 
        p_wishbone_bd_ram_mem3_111_31, p_wishbone_bd_ram_mem3_112_24, 
        p_wishbone_bd_ram_mem3_112_25, p_wishbone_bd_ram_mem3_112_26, 
        p_wishbone_bd_ram_mem3_112_27, p_wishbone_bd_ram_mem3_112_28, 
        p_wishbone_bd_ram_mem3_112_29, p_wishbone_bd_ram_mem3_112_30, 
        p_wishbone_bd_ram_mem3_112_31, p_wishbone_bd_ram_mem3_113_24, 
        p_wishbone_bd_ram_mem3_113_25, p_wishbone_bd_ram_mem3_113_26, 
        p_wishbone_bd_ram_mem3_113_27, p_wishbone_bd_ram_mem3_113_28, 
        p_wishbone_bd_ram_mem3_113_29, p_wishbone_bd_ram_mem3_113_30, 
        p_wishbone_bd_ram_mem3_113_31, p_wishbone_bd_ram_mem3_114_24, 
        p_wishbone_bd_ram_mem3_114_25, p_wishbone_bd_ram_mem3_114_26, 
        p_wishbone_bd_ram_mem3_114_27, p_wishbone_bd_ram_mem3_114_28, 
        p_wishbone_bd_ram_mem3_114_29, p_wishbone_bd_ram_mem3_114_30, 
        p_wishbone_bd_ram_mem3_114_31, p_wishbone_bd_ram_mem3_115_24, 
        p_wishbone_bd_ram_mem3_115_25, p_wishbone_bd_ram_mem3_115_26, 
        p_wishbone_bd_ram_mem3_115_27, p_wishbone_bd_ram_mem3_115_28, 
        p_wishbone_bd_ram_mem3_115_29, p_wishbone_bd_ram_mem3_115_30, 
        p_wishbone_bd_ram_mem3_115_31, p_wishbone_bd_ram_mem3_116_24, 
        p_wishbone_bd_ram_mem3_116_25, p_wishbone_bd_ram_mem3_116_26, 
        p_wishbone_bd_ram_mem3_116_27, p_wishbone_bd_ram_mem3_116_28, 
        p_wishbone_bd_ram_mem3_116_29, p_wishbone_bd_ram_mem3_116_30, 
        p_wishbone_bd_ram_mem3_116_31, p_wishbone_bd_ram_mem3_117_24, 
        p_wishbone_bd_ram_mem3_117_25, p_wishbone_bd_ram_mem3_117_26, 
        p_wishbone_bd_ram_mem3_117_27, p_wishbone_bd_ram_mem3_117_28, 
        p_wishbone_bd_ram_mem3_117_29, p_wishbone_bd_ram_mem3_117_30, 
        p_wishbone_bd_ram_mem3_117_31, p_wishbone_bd_ram_mem3_118_24, 
        p_wishbone_bd_ram_mem3_118_25, p_wishbone_bd_ram_mem3_118_26, 
        p_wishbone_bd_ram_mem3_118_27, p_wishbone_bd_ram_mem3_118_28, 
        p_wishbone_bd_ram_mem3_118_29, p_wishbone_bd_ram_mem3_118_30, 
        p_wishbone_bd_ram_mem3_118_31, p_wishbone_bd_ram_mem3_119_24, 
        p_wishbone_bd_ram_mem3_119_25, p_wishbone_bd_ram_mem3_119_26, 
        p_wishbone_bd_ram_mem3_119_27, p_wishbone_bd_ram_mem3_119_28, 
        p_wishbone_bd_ram_mem3_119_29, p_wishbone_bd_ram_mem3_119_30, 
        p_wishbone_bd_ram_mem3_119_31, p_wishbone_bd_ram_mem3_120_24, 
        p_wishbone_bd_ram_mem3_120_25, p_wishbone_bd_ram_mem3_120_26, 
        p_wishbone_bd_ram_mem3_120_27, p_wishbone_bd_ram_mem3_120_28, 
        p_wishbone_bd_ram_mem3_120_29, p_wishbone_bd_ram_mem3_120_30, 
        p_wishbone_bd_ram_mem3_120_31, p_wishbone_bd_ram_mem3_121_24, 
        p_wishbone_bd_ram_mem3_121_25, p_wishbone_bd_ram_mem3_121_26, 
        p_wishbone_bd_ram_mem3_121_27, p_wishbone_bd_ram_mem3_121_28, 
        p_wishbone_bd_ram_mem3_121_29, p_wishbone_bd_ram_mem3_121_30, 
        p_wishbone_bd_ram_mem3_121_31, p_wishbone_bd_ram_mem3_122_24, 
        p_wishbone_bd_ram_mem3_122_25, p_wishbone_bd_ram_mem3_122_26, 
        p_wishbone_bd_ram_mem3_122_27, p_wishbone_bd_ram_mem3_122_28, 
        p_wishbone_bd_ram_mem3_122_29, p_wishbone_bd_ram_mem3_122_30, 
        p_wishbone_bd_ram_mem3_122_31, p_wishbone_bd_ram_mem3_123_24, 
        p_wishbone_bd_ram_mem3_123_25, p_wishbone_bd_ram_mem3_123_26, 
        p_wishbone_bd_ram_mem3_123_27, p_wishbone_bd_ram_mem3_123_28, 
        p_wishbone_bd_ram_mem3_123_29, p_wishbone_bd_ram_mem3_123_30, 
        p_wishbone_bd_ram_mem3_123_31, p_wishbone_bd_ram_mem3_124_24, 
        p_wishbone_bd_ram_mem3_124_25, p_wishbone_bd_ram_mem3_124_26, 
        p_wishbone_bd_ram_mem3_124_27, p_wishbone_bd_ram_mem3_124_28, 
        p_wishbone_bd_ram_mem3_124_29, p_wishbone_bd_ram_mem3_124_30, 
        p_wishbone_bd_ram_mem3_124_31, p_wishbone_bd_ram_mem3_125_24, 
        p_wishbone_bd_ram_mem3_125_25, p_wishbone_bd_ram_mem3_125_26, 
        p_wishbone_bd_ram_mem3_125_27, p_wishbone_bd_ram_mem3_125_28, 
        p_wishbone_bd_ram_mem3_125_29, p_wishbone_bd_ram_mem3_125_30, 
        p_wishbone_bd_ram_mem3_125_31, p_wishbone_bd_ram_mem3_126_24, 
        p_wishbone_bd_ram_mem3_126_25, p_wishbone_bd_ram_mem3_126_26, 
        p_wishbone_bd_ram_mem3_126_27, p_wishbone_bd_ram_mem3_126_28, 
        p_wishbone_bd_ram_mem3_126_29, p_wishbone_bd_ram_mem3_126_30, 
        p_wishbone_bd_ram_mem3_126_31, p_wishbone_bd_ram_mem3_127_24, 
        p_wishbone_bd_ram_mem3_127_25, p_wishbone_bd_ram_mem3_127_26, 
        p_wishbone_bd_ram_mem3_127_27, p_wishbone_bd_ram_mem3_127_28, 
        p_wishbone_bd_ram_mem3_127_29, p_wishbone_bd_ram_mem3_127_30, 
        p_wishbone_bd_ram_mem3_127_31, p_wishbone_bd_ram_mem3_128_24, 
        p_wishbone_bd_ram_mem3_128_25, p_wishbone_bd_ram_mem3_128_26, 
        p_wishbone_bd_ram_mem3_128_27, p_wishbone_bd_ram_mem3_128_28, 
        p_wishbone_bd_ram_mem3_128_29, p_wishbone_bd_ram_mem3_128_30, 
        p_wishbone_bd_ram_mem3_128_31, p_wishbone_bd_ram_mem3_129_24, 
        p_wishbone_bd_ram_mem3_129_25, p_wishbone_bd_ram_mem3_129_26, 
        p_wishbone_bd_ram_mem3_129_27, p_wishbone_bd_ram_mem3_129_28, 
        p_wishbone_bd_ram_mem3_129_29, p_wishbone_bd_ram_mem3_129_30, 
        p_wishbone_bd_ram_mem3_129_31, p_wishbone_bd_ram_mem3_130_24, 
        p_wishbone_bd_ram_mem3_130_25, p_wishbone_bd_ram_mem3_130_26, 
        p_wishbone_bd_ram_mem3_130_27, p_wishbone_bd_ram_mem3_130_28, 
        p_wishbone_bd_ram_mem3_130_29, p_wishbone_bd_ram_mem3_130_30, 
        p_wishbone_bd_ram_mem3_130_31, p_wishbone_bd_ram_mem3_131_24, 
        p_wishbone_bd_ram_mem3_131_25, p_wishbone_bd_ram_mem3_131_26, 
        p_wishbone_bd_ram_mem3_131_27, p_wishbone_bd_ram_mem3_131_28, 
        p_wishbone_bd_ram_mem3_131_29, p_wishbone_bd_ram_mem3_131_30, 
        p_wishbone_bd_ram_mem3_131_31, p_wishbone_bd_ram_mem3_132_24, 
        p_wishbone_bd_ram_mem3_132_25, p_wishbone_bd_ram_mem3_132_26, 
        p_wishbone_bd_ram_mem3_132_27, p_wishbone_bd_ram_mem3_132_28, 
        p_wishbone_bd_ram_mem3_132_29, p_wishbone_bd_ram_mem3_132_30, 
        p_wishbone_bd_ram_mem3_132_31, p_wishbone_bd_ram_mem3_133_24, 
        p_wishbone_bd_ram_mem3_133_25, p_wishbone_bd_ram_mem3_133_26, 
        p_wishbone_bd_ram_mem3_133_27, p_wishbone_bd_ram_mem3_133_28, 
        p_wishbone_bd_ram_mem3_133_29, p_wishbone_bd_ram_mem3_133_30, 
        p_wishbone_bd_ram_mem3_133_31, p_wishbone_bd_ram_mem3_134_24, 
        p_wishbone_bd_ram_mem3_134_25, p_wishbone_bd_ram_mem3_134_26, 
        p_wishbone_bd_ram_mem3_134_27, p_wishbone_bd_ram_mem3_134_28, 
        p_wishbone_bd_ram_mem3_134_29, p_wishbone_bd_ram_mem3_134_30, 
        p_wishbone_bd_ram_mem3_134_31, p_wishbone_bd_ram_mem3_135_24, 
        p_wishbone_bd_ram_mem3_135_25, p_wishbone_bd_ram_mem3_135_26, 
        p_wishbone_bd_ram_mem3_135_27, p_wishbone_bd_ram_mem3_135_28, 
        p_wishbone_bd_ram_mem3_135_29, p_wishbone_bd_ram_mem3_135_30, 
        p_wishbone_bd_ram_mem3_135_31, p_wishbone_bd_ram_mem3_136_24, 
        p_wishbone_bd_ram_mem3_136_25, p_wishbone_bd_ram_mem3_136_26, 
        p_wishbone_bd_ram_mem3_136_27, p_wishbone_bd_ram_mem3_136_28, 
        p_wishbone_bd_ram_mem3_136_29, p_wishbone_bd_ram_mem3_136_30, 
        p_wishbone_bd_ram_mem3_136_31, p_wishbone_bd_ram_mem3_137_24, 
        p_wishbone_bd_ram_mem3_137_25, p_wishbone_bd_ram_mem3_137_26, 
        p_wishbone_bd_ram_mem3_137_27, p_wishbone_bd_ram_mem3_137_28, 
        p_wishbone_bd_ram_mem3_137_29, p_wishbone_bd_ram_mem3_137_30, 
        p_wishbone_bd_ram_mem3_137_31, p_wishbone_bd_ram_mem3_138_24, 
        p_wishbone_bd_ram_mem3_138_25, p_wishbone_bd_ram_mem3_138_26, 
        p_wishbone_bd_ram_mem3_138_27, p_wishbone_bd_ram_mem3_138_28, 
        p_wishbone_bd_ram_mem3_138_29, p_wishbone_bd_ram_mem3_138_30, 
        p_wishbone_bd_ram_mem3_138_31, p_wishbone_bd_ram_mem3_139_24, 
        p_wishbone_bd_ram_mem3_139_25, p_wishbone_bd_ram_mem3_139_26, 
        p_wishbone_bd_ram_mem3_139_27, p_wishbone_bd_ram_mem3_139_28, 
        p_wishbone_bd_ram_mem3_139_29, p_wishbone_bd_ram_mem3_139_30, 
        p_wishbone_bd_ram_mem3_139_31, p_wishbone_bd_ram_mem3_140_24, 
        p_wishbone_bd_ram_mem3_140_25, p_wishbone_bd_ram_mem3_140_26, 
        p_wishbone_bd_ram_mem3_140_27, p_wishbone_bd_ram_mem3_140_28, 
        p_wishbone_bd_ram_mem3_140_29, p_wishbone_bd_ram_mem3_140_30, 
        p_wishbone_bd_ram_mem3_140_31, p_wishbone_bd_ram_mem3_141_24, 
        p_wishbone_bd_ram_mem3_141_25, p_wishbone_bd_ram_mem3_141_26, 
        p_wishbone_bd_ram_mem3_141_27, p_wishbone_bd_ram_mem3_141_28, 
        p_wishbone_bd_ram_mem3_141_29, p_wishbone_bd_ram_mem3_141_30, 
        p_wishbone_bd_ram_mem3_141_31, p_wishbone_bd_ram_mem3_142_24, 
        p_wishbone_bd_ram_mem3_142_25, p_wishbone_bd_ram_mem3_142_26, 
        p_wishbone_bd_ram_mem3_142_27, p_wishbone_bd_ram_mem3_142_28, 
        p_wishbone_bd_ram_mem3_142_29, p_wishbone_bd_ram_mem3_142_30, 
        p_wishbone_bd_ram_mem3_142_31, p_wishbone_bd_ram_mem3_143_24, 
        p_wishbone_bd_ram_mem3_143_25, p_wishbone_bd_ram_mem3_143_26, 
        p_wishbone_bd_ram_mem3_143_27, p_wishbone_bd_ram_mem3_143_28, 
        p_wishbone_bd_ram_mem3_143_29, p_wishbone_bd_ram_mem3_143_30, 
        p_wishbone_bd_ram_mem3_143_31, p_wishbone_bd_ram_mem3_144_24, 
        p_wishbone_bd_ram_mem3_144_25, p_wishbone_bd_ram_mem3_144_26, 
        p_wishbone_bd_ram_mem3_144_27, p_wishbone_bd_ram_mem3_144_28, 
        p_wishbone_bd_ram_mem3_144_29, p_wishbone_bd_ram_mem3_144_30, 
        p_wishbone_bd_ram_mem3_144_31, p_wishbone_bd_ram_mem3_145_24, 
        p_wishbone_bd_ram_mem3_145_25, p_wishbone_bd_ram_mem3_145_26, 
        p_wishbone_bd_ram_mem3_145_27, p_wishbone_bd_ram_mem3_145_28, 
        p_wishbone_bd_ram_mem3_145_29, p_wishbone_bd_ram_mem3_145_30, 
        p_wishbone_bd_ram_mem3_145_31, p_wishbone_bd_ram_mem3_146_24, 
        p_wishbone_bd_ram_mem3_146_25, p_wishbone_bd_ram_mem3_146_26, 
        p_wishbone_bd_ram_mem3_146_27, p_wishbone_bd_ram_mem3_146_28, 
        p_wishbone_bd_ram_mem3_146_29, p_wishbone_bd_ram_mem3_146_30, 
        p_wishbone_bd_ram_mem3_146_31, p_wishbone_bd_ram_mem3_147_24, 
        p_wishbone_bd_ram_mem3_147_25, p_wishbone_bd_ram_mem3_147_26, 
        p_wishbone_bd_ram_mem3_147_27, p_wishbone_bd_ram_mem3_147_28, 
        p_wishbone_bd_ram_mem3_147_29, p_wishbone_bd_ram_mem3_147_30, 
        p_wishbone_bd_ram_mem3_147_31, p_wishbone_bd_ram_mem3_148_24, 
        p_wishbone_bd_ram_mem3_148_25, p_wishbone_bd_ram_mem3_148_26, 
        p_wishbone_bd_ram_mem3_148_27, p_wishbone_bd_ram_mem3_148_28, 
        p_wishbone_bd_ram_mem3_148_29, p_wishbone_bd_ram_mem3_148_30, 
        p_wishbone_bd_ram_mem3_148_31, p_wishbone_bd_ram_mem3_149_24, 
        p_wishbone_bd_ram_mem3_149_25, p_wishbone_bd_ram_mem3_149_26, 
        p_wishbone_bd_ram_mem3_149_27, p_wishbone_bd_ram_mem3_149_28, 
        p_wishbone_bd_ram_mem3_149_29, p_wishbone_bd_ram_mem3_149_30, 
        p_wishbone_bd_ram_mem3_149_31, p_wishbone_bd_ram_mem3_150_24, 
        p_wishbone_bd_ram_mem3_150_25, p_wishbone_bd_ram_mem3_150_26, 
        p_wishbone_bd_ram_mem3_150_27, p_wishbone_bd_ram_mem3_150_28, 
        p_wishbone_bd_ram_mem3_150_29, p_wishbone_bd_ram_mem3_150_30, 
        p_wishbone_bd_ram_mem3_150_31, p_wishbone_bd_ram_mem3_151_24, 
        p_wishbone_bd_ram_mem3_151_25, p_wishbone_bd_ram_mem3_151_26, 
        p_wishbone_bd_ram_mem3_151_27, p_wishbone_bd_ram_mem3_151_28, 
        p_wishbone_bd_ram_mem3_151_29, p_wishbone_bd_ram_mem3_151_30, 
        p_wishbone_bd_ram_mem3_151_31, p_wishbone_bd_ram_mem3_152_24, 
        p_wishbone_bd_ram_mem3_152_25, p_wishbone_bd_ram_mem3_152_26, 
        p_wishbone_bd_ram_mem3_152_27, p_wishbone_bd_ram_mem3_152_28, 
        p_wishbone_bd_ram_mem3_152_29, p_wishbone_bd_ram_mem3_152_30, 
        p_wishbone_bd_ram_mem3_152_31, p_wishbone_bd_ram_mem3_153_24, 
        p_wishbone_bd_ram_mem3_153_25, p_wishbone_bd_ram_mem3_153_26, 
        p_wishbone_bd_ram_mem3_153_27, p_wishbone_bd_ram_mem3_153_28, 
        p_wishbone_bd_ram_mem3_153_29, p_wishbone_bd_ram_mem3_153_30, 
        p_wishbone_bd_ram_mem3_153_31, p_wishbone_bd_ram_mem3_154_24, 
        p_wishbone_bd_ram_mem3_154_25, p_wishbone_bd_ram_mem3_154_26, 
        p_wishbone_bd_ram_mem3_154_27, p_wishbone_bd_ram_mem3_154_28, 
        p_wishbone_bd_ram_mem3_154_29, p_wishbone_bd_ram_mem3_154_30, 
        p_wishbone_bd_ram_mem3_154_31, p_wishbone_bd_ram_mem3_155_24, 
        p_wishbone_bd_ram_mem3_155_25, p_wishbone_bd_ram_mem3_155_26, 
        p_wishbone_bd_ram_mem3_155_27, p_wishbone_bd_ram_mem3_155_28, 
        p_wishbone_bd_ram_mem3_155_29, p_wishbone_bd_ram_mem3_155_30, 
        p_wishbone_bd_ram_mem3_155_31, p_wishbone_bd_ram_mem3_156_24, 
        p_wishbone_bd_ram_mem3_156_25, p_wishbone_bd_ram_mem3_156_26, 
        p_wishbone_bd_ram_mem3_156_27, p_wishbone_bd_ram_mem3_156_28, 
        p_wishbone_bd_ram_mem3_156_29, p_wishbone_bd_ram_mem3_156_30, 
        p_wishbone_bd_ram_mem3_156_31, p_wishbone_bd_ram_mem3_157_24, 
        p_wishbone_bd_ram_mem3_157_25, p_wishbone_bd_ram_mem3_157_26, 
        p_wishbone_bd_ram_mem3_157_27, p_wishbone_bd_ram_mem3_157_28, 
        p_wishbone_bd_ram_mem3_157_29, p_wishbone_bd_ram_mem3_157_30, 
        p_wishbone_bd_ram_mem3_157_31, p_wishbone_bd_ram_mem3_158_24, 
        p_wishbone_bd_ram_mem3_158_25, p_wishbone_bd_ram_mem3_158_26, 
        p_wishbone_bd_ram_mem3_158_27, p_wishbone_bd_ram_mem3_158_28, 
        p_wishbone_bd_ram_mem3_158_29, p_wishbone_bd_ram_mem3_158_30, 
        p_wishbone_bd_ram_mem3_158_31, p_wishbone_bd_ram_mem3_159_24, 
        p_wishbone_bd_ram_mem3_159_25, p_wishbone_bd_ram_mem3_159_26, 
        p_wishbone_bd_ram_mem3_159_27, p_wishbone_bd_ram_mem3_159_28, 
        p_wishbone_bd_ram_mem3_159_29, p_wishbone_bd_ram_mem3_159_30, 
        p_wishbone_bd_ram_mem3_159_31, p_wishbone_bd_ram_mem3_160_24, 
        p_wishbone_bd_ram_mem3_160_25, p_wishbone_bd_ram_mem3_160_26, 
        p_wishbone_bd_ram_mem3_160_27, p_wishbone_bd_ram_mem3_160_28, 
        p_wishbone_bd_ram_mem3_160_29, p_wishbone_bd_ram_mem3_160_30, 
        p_wishbone_bd_ram_mem3_160_31, p_wishbone_bd_ram_mem3_161_24, 
        p_wishbone_bd_ram_mem3_161_25, p_wishbone_bd_ram_mem3_161_26, 
        p_wishbone_bd_ram_mem3_161_27, p_wishbone_bd_ram_mem3_161_28, 
        p_wishbone_bd_ram_mem3_161_29, p_wishbone_bd_ram_mem3_161_30, 
        p_wishbone_bd_ram_mem3_161_31, p_wishbone_bd_ram_mem3_162_24, 
        p_wishbone_bd_ram_mem3_162_25, p_wishbone_bd_ram_mem3_162_26, 
        p_wishbone_bd_ram_mem3_162_27, p_wishbone_bd_ram_mem3_162_28, 
        p_wishbone_bd_ram_mem3_162_29, p_wishbone_bd_ram_mem3_162_30, 
        p_wishbone_bd_ram_mem3_162_31, p_wishbone_bd_ram_mem3_163_24, 
        p_wishbone_bd_ram_mem3_163_25, p_wishbone_bd_ram_mem3_163_26, 
        p_wishbone_bd_ram_mem3_163_27, p_wishbone_bd_ram_mem3_163_28, 
        p_wishbone_bd_ram_mem3_163_29, p_wishbone_bd_ram_mem3_163_30, 
        p_wishbone_bd_ram_mem3_163_31, p_wishbone_bd_ram_mem3_164_24, 
        p_wishbone_bd_ram_mem3_164_25, p_wishbone_bd_ram_mem3_164_26, 
        p_wishbone_bd_ram_mem3_164_27, p_wishbone_bd_ram_mem3_164_28, 
        p_wishbone_bd_ram_mem3_164_29, p_wishbone_bd_ram_mem3_164_30, 
        p_wishbone_bd_ram_mem3_164_31, p_wishbone_bd_ram_mem3_165_24, 
        p_wishbone_bd_ram_mem3_165_25, p_wishbone_bd_ram_mem3_165_26, 
        p_wishbone_bd_ram_mem3_165_27, p_wishbone_bd_ram_mem3_165_28, 
        p_wishbone_bd_ram_mem3_165_29, p_wishbone_bd_ram_mem3_165_30, 
        p_wishbone_bd_ram_mem3_165_31, p_wishbone_bd_ram_mem3_166_24, 
        p_wishbone_bd_ram_mem3_166_25, p_wishbone_bd_ram_mem3_166_26, 
        p_wishbone_bd_ram_mem3_166_27, p_wishbone_bd_ram_mem3_166_28, 
        p_wishbone_bd_ram_mem3_166_29, p_wishbone_bd_ram_mem3_166_30, 
        p_wishbone_bd_ram_mem3_166_31, p_wishbone_bd_ram_mem3_167_24, 
        p_wishbone_bd_ram_mem3_167_25, p_wishbone_bd_ram_mem3_167_26, 
        p_wishbone_bd_ram_mem3_167_27, p_wishbone_bd_ram_mem3_167_28, 
        p_wishbone_bd_ram_mem3_167_29, p_wishbone_bd_ram_mem3_167_30, 
        p_wishbone_bd_ram_mem3_167_31, p_wishbone_bd_ram_mem3_168_24, 
        p_wishbone_bd_ram_mem3_168_25, p_wishbone_bd_ram_mem3_168_26, 
        p_wishbone_bd_ram_mem3_168_27, p_wishbone_bd_ram_mem3_168_28, 
        p_wishbone_bd_ram_mem3_168_29, p_wishbone_bd_ram_mem3_168_30, 
        p_wishbone_bd_ram_mem3_168_31, p_wishbone_bd_ram_mem3_169_24, 
        p_wishbone_bd_ram_mem3_169_25, p_wishbone_bd_ram_mem3_169_26, 
        p_wishbone_bd_ram_mem3_169_27, p_wishbone_bd_ram_mem3_169_28, 
        p_wishbone_bd_ram_mem3_169_29, p_wishbone_bd_ram_mem3_169_30, 
        p_wishbone_bd_ram_mem3_169_31, p_wishbone_bd_ram_mem3_170_24, 
        p_wishbone_bd_ram_mem3_170_25, p_wishbone_bd_ram_mem3_170_26, 
        p_wishbone_bd_ram_mem3_170_27, p_wishbone_bd_ram_mem3_170_28, 
        p_wishbone_bd_ram_mem3_170_29, p_wishbone_bd_ram_mem3_170_30, 
        p_wishbone_bd_ram_mem3_170_31, p_wishbone_bd_ram_mem3_171_24, 
        p_wishbone_bd_ram_mem3_171_25, p_wishbone_bd_ram_mem3_171_26, 
        p_wishbone_bd_ram_mem3_171_27, p_wishbone_bd_ram_mem3_171_28, 
        p_wishbone_bd_ram_mem3_171_29, p_wishbone_bd_ram_mem3_171_30, 
        p_wishbone_bd_ram_mem3_171_31, p_wishbone_bd_ram_mem3_172_24, 
        p_wishbone_bd_ram_mem3_172_25, p_wishbone_bd_ram_mem3_172_26, 
        p_wishbone_bd_ram_mem3_172_27, p_wishbone_bd_ram_mem3_172_28, 
        p_wishbone_bd_ram_mem3_172_29, p_wishbone_bd_ram_mem3_172_30, 
        p_wishbone_bd_ram_mem3_172_31, p_wishbone_bd_ram_mem3_173_24, 
        p_wishbone_bd_ram_mem3_173_25, p_wishbone_bd_ram_mem3_173_26, 
        p_wishbone_bd_ram_mem3_173_27, p_wishbone_bd_ram_mem3_173_28, 
        p_wishbone_bd_ram_mem3_173_29, p_wishbone_bd_ram_mem3_173_30, 
        p_wishbone_bd_ram_mem3_173_31, p_wishbone_bd_ram_mem3_174_24, 
        p_wishbone_bd_ram_mem3_174_25, p_wishbone_bd_ram_mem3_174_26, 
        p_wishbone_bd_ram_mem3_174_27, p_wishbone_bd_ram_mem3_174_28, 
        p_wishbone_bd_ram_mem3_174_29, p_wishbone_bd_ram_mem3_174_30, 
        p_wishbone_bd_ram_mem3_174_31, p_wishbone_bd_ram_mem3_175_24, 
        p_wishbone_bd_ram_mem3_175_25, p_wishbone_bd_ram_mem3_175_26, 
        p_wishbone_bd_ram_mem3_175_27, p_wishbone_bd_ram_mem3_175_28, 
        p_wishbone_bd_ram_mem3_175_29, p_wishbone_bd_ram_mem3_175_30, 
        p_wishbone_bd_ram_mem3_175_31, p_wishbone_bd_ram_mem3_176_24, 
        p_wishbone_bd_ram_mem3_176_25, p_wishbone_bd_ram_mem3_176_26, 
        p_wishbone_bd_ram_mem3_176_27, p_wishbone_bd_ram_mem3_176_28, 
        p_wishbone_bd_ram_mem3_176_29, p_wishbone_bd_ram_mem3_176_30, 
        p_wishbone_bd_ram_mem3_176_31, p_wishbone_bd_ram_mem3_177_24, 
        p_wishbone_bd_ram_mem3_177_25, p_wishbone_bd_ram_mem3_177_26, 
        p_wishbone_bd_ram_mem3_177_27, p_wishbone_bd_ram_mem3_177_28, 
        p_wishbone_bd_ram_mem3_177_29, p_wishbone_bd_ram_mem3_177_30, 
        p_wishbone_bd_ram_mem3_177_31, p_wishbone_bd_ram_mem3_178_24, 
        p_wishbone_bd_ram_mem3_178_25, p_wishbone_bd_ram_mem3_178_26, 
        p_wishbone_bd_ram_mem3_178_27, p_wishbone_bd_ram_mem3_178_28, 
        p_wishbone_bd_ram_mem3_178_29, p_wishbone_bd_ram_mem3_178_30, 
        p_wishbone_bd_ram_mem3_178_31, p_wishbone_bd_ram_mem3_179_24, 
        p_wishbone_bd_ram_mem3_179_25, p_wishbone_bd_ram_mem3_179_26, 
        p_wishbone_bd_ram_mem3_179_27, p_wishbone_bd_ram_mem3_179_28, 
        p_wishbone_bd_ram_mem3_179_29, p_wishbone_bd_ram_mem3_179_30, 
        p_wishbone_bd_ram_mem3_179_31, p_wishbone_bd_ram_mem3_180_24, 
        p_wishbone_bd_ram_mem3_180_25, p_wishbone_bd_ram_mem3_180_26, 
        p_wishbone_bd_ram_mem3_180_27, p_wishbone_bd_ram_mem3_180_28, 
        p_wishbone_bd_ram_mem3_180_29, p_wishbone_bd_ram_mem3_180_30, 
        p_wishbone_bd_ram_mem3_180_31, p_wishbone_bd_ram_mem3_181_24, 
        p_wishbone_bd_ram_mem3_181_25, p_wishbone_bd_ram_mem3_181_26, 
        p_wishbone_bd_ram_mem3_181_27, p_wishbone_bd_ram_mem3_181_28, 
        p_wishbone_bd_ram_mem3_181_29, p_wishbone_bd_ram_mem3_181_30, 
        p_wishbone_bd_ram_mem3_181_31, p_wishbone_bd_ram_mem3_182_24, 
        p_wishbone_bd_ram_mem3_182_25, p_wishbone_bd_ram_mem3_182_26, 
        p_wishbone_bd_ram_mem3_182_27, p_wishbone_bd_ram_mem3_182_28, 
        p_wishbone_bd_ram_mem3_182_29, p_wishbone_bd_ram_mem3_182_30, 
        p_wishbone_bd_ram_mem3_182_31, p_wishbone_bd_ram_mem3_183_24, 
        p_wishbone_bd_ram_mem3_183_25, p_wishbone_bd_ram_mem3_183_26, 
        p_wishbone_bd_ram_mem3_183_27, p_wishbone_bd_ram_mem3_183_28, 
        p_wishbone_bd_ram_mem3_183_29, p_wishbone_bd_ram_mem3_183_30, 
        p_wishbone_bd_ram_mem3_183_31, p_wishbone_bd_ram_mem3_184_24, 
        p_wishbone_bd_ram_mem3_184_25, p_wishbone_bd_ram_mem3_184_26, 
        p_wishbone_bd_ram_mem3_184_27, p_wishbone_bd_ram_mem3_184_28, 
        p_wishbone_bd_ram_mem3_184_29, p_wishbone_bd_ram_mem3_184_30, 
        p_wishbone_bd_ram_mem3_184_31, p_wishbone_bd_ram_mem3_185_24, 
        p_wishbone_bd_ram_mem3_185_25, p_wishbone_bd_ram_mem3_185_26, 
        p_wishbone_bd_ram_mem3_185_27, p_wishbone_bd_ram_mem3_185_28, 
        p_wishbone_bd_ram_mem3_185_29, p_wishbone_bd_ram_mem3_185_30, 
        p_wishbone_bd_ram_mem3_185_31, p_wishbone_bd_ram_mem3_186_24, 
        p_wishbone_bd_ram_mem3_186_25, p_wishbone_bd_ram_mem3_186_26, 
        p_wishbone_bd_ram_mem3_186_27, p_wishbone_bd_ram_mem3_186_28, 
        p_wishbone_bd_ram_mem3_186_29, p_wishbone_bd_ram_mem3_186_30, 
        p_wishbone_bd_ram_mem3_186_31, p_wishbone_bd_ram_mem3_187_24, 
        p_wishbone_bd_ram_mem3_187_25, p_wishbone_bd_ram_mem3_187_26, 
        p_wishbone_bd_ram_mem3_187_27, p_wishbone_bd_ram_mem3_187_28, 
        p_wishbone_bd_ram_mem3_187_29, p_wishbone_bd_ram_mem3_187_30, 
        p_wishbone_bd_ram_mem3_187_31, p_wishbone_bd_ram_mem3_188_24, 
        p_wishbone_bd_ram_mem3_188_25, p_wishbone_bd_ram_mem3_188_26, 
        p_wishbone_bd_ram_mem3_188_27, p_wishbone_bd_ram_mem3_188_28, 
        p_wishbone_bd_ram_mem3_188_29, p_wishbone_bd_ram_mem3_188_30, 
        p_wishbone_bd_ram_mem3_188_31, p_wishbone_bd_ram_mem3_189_24, 
        p_wishbone_bd_ram_mem3_189_25, p_wishbone_bd_ram_mem3_189_26, 
        p_wishbone_bd_ram_mem3_189_27, p_wishbone_bd_ram_mem3_189_28, 
        p_wishbone_bd_ram_mem3_189_29, p_wishbone_bd_ram_mem3_189_30, 
        p_wishbone_bd_ram_mem3_189_31, p_wishbone_bd_ram_mem3_190_24, 
        p_wishbone_bd_ram_mem3_190_25, p_wishbone_bd_ram_mem3_190_26, 
        p_wishbone_bd_ram_mem3_190_27, p_wishbone_bd_ram_mem3_190_28, 
        p_wishbone_bd_ram_mem3_190_29, p_wishbone_bd_ram_mem3_190_30, 
        p_wishbone_bd_ram_mem3_190_31, p_wishbone_bd_ram_mem3_191_24, 
        p_wishbone_bd_ram_mem3_191_25, p_wishbone_bd_ram_mem3_191_26, 
        p_wishbone_bd_ram_mem3_191_27, p_wishbone_bd_ram_mem3_191_28, 
        p_wishbone_bd_ram_mem3_191_29, p_wishbone_bd_ram_mem3_191_30, 
        p_wishbone_bd_ram_mem3_191_31, p_wishbone_bd_ram_mem3_192_24, 
        p_wishbone_bd_ram_mem3_192_25, p_wishbone_bd_ram_mem3_192_26, 
        p_wishbone_bd_ram_mem3_192_27, p_wishbone_bd_ram_mem3_192_28, 
        p_wishbone_bd_ram_mem3_192_29, p_wishbone_bd_ram_mem3_192_30, 
        p_wishbone_bd_ram_mem3_192_31, p_wishbone_bd_ram_mem3_193_24, 
        p_wishbone_bd_ram_mem3_193_25, p_wishbone_bd_ram_mem3_193_26, 
        p_wishbone_bd_ram_mem3_193_27, p_wishbone_bd_ram_mem3_193_28, 
        p_wishbone_bd_ram_mem3_193_29, p_wishbone_bd_ram_mem3_193_30, 
        p_wishbone_bd_ram_mem3_193_31, p_wishbone_bd_ram_mem3_194_24, 
        p_wishbone_bd_ram_mem3_194_25, p_wishbone_bd_ram_mem3_194_26, 
        p_wishbone_bd_ram_mem3_194_27, p_wishbone_bd_ram_mem3_194_28, 
        p_wishbone_bd_ram_mem3_194_29, p_wishbone_bd_ram_mem3_194_30, 
        p_wishbone_bd_ram_mem3_194_31, p_wishbone_bd_ram_mem3_195_24, 
        p_wishbone_bd_ram_mem3_195_25, p_wishbone_bd_ram_mem3_195_26, 
        p_wishbone_bd_ram_mem3_195_27, p_wishbone_bd_ram_mem3_195_28, 
        p_wishbone_bd_ram_mem3_195_29, p_wishbone_bd_ram_mem3_195_30, 
        p_wishbone_bd_ram_mem3_195_31, p_wishbone_bd_ram_mem3_196_24, 
        p_wishbone_bd_ram_mem3_196_25, p_wishbone_bd_ram_mem3_196_26, 
        p_wishbone_bd_ram_mem3_196_27, p_wishbone_bd_ram_mem3_196_28, 
        p_wishbone_bd_ram_mem3_196_29, p_wishbone_bd_ram_mem3_196_30, 
        p_wishbone_bd_ram_mem3_196_31, p_wishbone_bd_ram_mem3_197_24, 
        p_wishbone_bd_ram_mem3_197_25, p_wishbone_bd_ram_mem3_197_26, 
        p_wishbone_bd_ram_mem3_197_27, p_wishbone_bd_ram_mem3_197_28, 
        p_wishbone_bd_ram_mem3_197_29, p_wishbone_bd_ram_mem3_197_30, 
        p_wishbone_bd_ram_mem3_197_31, p_wishbone_bd_ram_mem3_198_24, 
        p_wishbone_bd_ram_mem3_198_25, p_wishbone_bd_ram_mem3_198_26, 
        p_wishbone_bd_ram_mem3_198_27, p_wishbone_bd_ram_mem3_198_28, 
        p_wishbone_bd_ram_mem3_198_29, p_wishbone_bd_ram_mem3_198_30, 
        p_wishbone_bd_ram_mem3_198_31, p_wishbone_bd_ram_mem3_199_24, 
        p_wishbone_bd_ram_mem3_199_25, p_wishbone_bd_ram_mem3_199_26, 
        p_wishbone_bd_ram_mem3_199_27, p_wishbone_bd_ram_mem3_199_28, 
        p_wishbone_bd_ram_mem3_199_29, p_wishbone_bd_ram_mem3_199_30, 
        p_wishbone_bd_ram_mem3_199_31, p_wishbone_bd_ram_mem3_200_24, 
        p_wishbone_bd_ram_mem3_200_25, p_wishbone_bd_ram_mem3_200_26, 
        p_wishbone_bd_ram_mem3_200_27, p_wishbone_bd_ram_mem3_200_28, 
        p_wishbone_bd_ram_mem3_200_29, p_wishbone_bd_ram_mem3_200_30, 
        p_wishbone_bd_ram_mem3_200_31, p_wishbone_bd_ram_mem3_201_24, 
        p_wishbone_bd_ram_mem3_201_25, p_wishbone_bd_ram_mem3_201_26, 
        p_wishbone_bd_ram_mem3_201_27, p_wishbone_bd_ram_mem3_201_28, 
        p_wishbone_bd_ram_mem3_201_29, p_wishbone_bd_ram_mem3_201_30, 
        p_wishbone_bd_ram_mem3_201_31, p_wishbone_bd_ram_mem3_202_24, 
        p_wishbone_bd_ram_mem3_202_25, p_wishbone_bd_ram_mem3_202_26, 
        p_wishbone_bd_ram_mem3_202_27, p_wishbone_bd_ram_mem3_202_28, 
        p_wishbone_bd_ram_mem3_202_29, p_wishbone_bd_ram_mem3_202_30, 
        p_wishbone_bd_ram_mem3_202_31, p_wishbone_bd_ram_mem3_203_24, 
        p_wishbone_bd_ram_mem3_203_25, p_wishbone_bd_ram_mem3_203_26, 
        p_wishbone_bd_ram_mem3_203_27, p_wishbone_bd_ram_mem3_203_28, 
        p_wishbone_bd_ram_mem3_203_29, p_wishbone_bd_ram_mem3_203_30, 
        p_wishbone_bd_ram_mem3_203_31, p_wishbone_bd_ram_mem3_204_24, 
        p_wishbone_bd_ram_mem3_204_25, p_wishbone_bd_ram_mem3_204_26, 
        p_wishbone_bd_ram_mem3_204_27, p_wishbone_bd_ram_mem3_204_28, 
        p_wishbone_bd_ram_mem3_204_29, p_wishbone_bd_ram_mem3_204_30, 
        p_wishbone_bd_ram_mem3_204_31, p_wishbone_bd_ram_mem3_205_24, 
        p_wishbone_bd_ram_mem3_205_25, p_wishbone_bd_ram_mem3_205_26, 
        p_wishbone_bd_ram_mem3_205_27, p_wishbone_bd_ram_mem3_205_28, 
        p_wishbone_bd_ram_mem3_205_29, p_wishbone_bd_ram_mem3_205_30, 
        p_wishbone_bd_ram_mem3_205_31, p_wishbone_bd_ram_mem3_206_24, 
        p_wishbone_bd_ram_mem3_206_25, p_wishbone_bd_ram_mem3_206_26, 
        p_wishbone_bd_ram_mem3_206_27, p_wishbone_bd_ram_mem3_206_28, 
        p_wishbone_bd_ram_mem3_206_29, p_wishbone_bd_ram_mem3_206_30, 
        p_wishbone_bd_ram_mem3_206_31, p_wishbone_bd_ram_mem3_207_24, 
        p_wishbone_bd_ram_mem3_207_25, p_wishbone_bd_ram_mem3_207_26, 
        p_wishbone_bd_ram_mem3_207_27, p_wishbone_bd_ram_mem3_207_28, 
        p_wishbone_bd_ram_mem3_207_29, p_wishbone_bd_ram_mem3_207_30, 
        p_wishbone_bd_ram_mem3_207_31, p_wishbone_bd_ram_mem3_208_24, 
        p_wishbone_bd_ram_mem3_208_25, p_wishbone_bd_ram_mem3_208_26, 
        p_wishbone_bd_ram_mem3_208_27, p_wishbone_bd_ram_mem3_208_28, 
        p_wishbone_bd_ram_mem3_208_29, p_wishbone_bd_ram_mem3_208_30, 
        p_wishbone_bd_ram_mem3_208_31, p_wishbone_bd_ram_mem3_209_24, 
        p_wishbone_bd_ram_mem3_209_25, p_wishbone_bd_ram_mem3_209_26, 
        p_wishbone_bd_ram_mem3_209_27, p_wishbone_bd_ram_mem3_209_28, 
        p_wishbone_bd_ram_mem3_209_29, p_wishbone_bd_ram_mem3_209_30, 
        p_wishbone_bd_ram_mem3_209_31, p_wishbone_bd_ram_mem3_210_24, 
        p_wishbone_bd_ram_mem3_210_25, p_wishbone_bd_ram_mem3_210_26, 
        p_wishbone_bd_ram_mem3_210_27, p_wishbone_bd_ram_mem3_210_28, 
        p_wishbone_bd_ram_mem3_210_29, p_wishbone_bd_ram_mem3_210_30, 
        p_wishbone_bd_ram_mem3_210_31, p_wishbone_bd_ram_mem3_211_24, 
        p_wishbone_bd_ram_mem3_211_25, p_wishbone_bd_ram_mem3_211_26, 
        p_wishbone_bd_ram_mem3_211_27, p_wishbone_bd_ram_mem3_211_28, 
        p_wishbone_bd_ram_mem3_211_29, p_wishbone_bd_ram_mem3_211_30, 
        p_wishbone_bd_ram_mem3_211_31, p_wishbone_bd_ram_mem3_212_24, 
        p_wishbone_bd_ram_mem3_212_25, p_wishbone_bd_ram_mem3_212_26, 
        p_wishbone_bd_ram_mem3_212_27, p_wishbone_bd_ram_mem3_212_28, 
        p_wishbone_bd_ram_mem3_212_29, p_wishbone_bd_ram_mem3_212_30, 
        p_wishbone_bd_ram_mem3_212_31, p_wishbone_bd_ram_mem3_213_24, 
        p_wishbone_bd_ram_mem3_213_25, p_wishbone_bd_ram_mem3_213_26, 
        p_wishbone_bd_ram_mem3_213_27, p_wishbone_bd_ram_mem3_213_28, 
        p_wishbone_bd_ram_mem3_213_29, p_wishbone_bd_ram_mem3_213_30, 
        p_wishbone_bd_ram_mem3_213_31, p_wishbone_bd_ram_mem3_214_24, 
        p_wishbone_bd_ram_mem3_214_25, p_wishbone_bd_ram_mem3_214_26, 
        p_wishbone_bd_ram_mem3_214_27, p_wishbone_bd_ram_mem3_214_28, 
        p_wishbone_bd_ram_mem3_214_29, p_wishbone_bd_ram_mem3_214_30, 
        p_wishbone_bd_ram_mem3_214_31, p_wishbone_bd_ram_mem3_215_24, 
        p_wishbone_bd_ram_mem3_215_25, p_wishbone_bd_ram_mem3_215_26, 
        p_wishbone_bd_ram_mem3_215_27, p_wishbone_bd_ram_mem3_215_28, 
        p_wishbone_bd_ram_mem3_215_29, p_wishbone_bd_ram_mem3_215_30, 
        p_wishbone_bd_ram_mem3_215_31, p_wishbone_bd_ram_mem3_216_24, 
        p_wishbone_bd_ram_mem3_216_25, p_wishbone_bd_ram_mem3_216_26, 
        p_wishbone_bd_ram_mem3_216_27, p_wishbone_bd_ram_mem3_216_28, 
        p_wishbone_bd_ram_mem3_216_29, p_wishbone_bd_ram_mem3_216_30, 
        p_wishbone_bd_ram_mem3_216_31, p_wishbone_bd_ram_mem3_217_24, 
        p_wishbone_bd_ram_mem3_217_25, p_wishbone_bd_ram_mem3_217_26, 
        p_wishbone_bd_ram_mem3_217_27, p_wishbone_bd_ram_mem3_217_28, 
        p_wishbone_bd_ram_mem3_217_29, p_wishbone_bd_ram_mem3_217_30, 
        p_wishbone_bd_ram_mem3_217_31, p_wishbone_bd_ram_mem3_218_24, 
        p_wishbone_bd_ram_mem3_218_25, p_wishbone_bd_ram_mem3_218_26, 
        p_wishbone_bd_ram_mem3_218_27, p_wishbone_bd_ram_mem3_218_28, 
        p_wishbone_bd_ram_mem3_218_29, p_wishbone_bd_ram_mem3_218_30, 
        p_wishbone_bd_ram_mem3_218_31, p_wishbone_bd_ram_mem3_219_24, 
        p_wishbone_bd_ram_mem3_219_25, p_wishbone_bd_ram_mem3_219_26, 
        p_wishbone_bd_ram_mem3_219_27, p_wishbone_bd_ram_mem3_219_28, 
        p_wishbone_bd_ram_mem3_219_29, p_wishbone_bd_ram_mem3_219_30, 
        p_wishbone_bd_ram_mem3_219_31, p_wishbone_bd_ram_mem3_220_24, 
        p_wishbone_bd_ram_mem3_220_25, p_wishbone_bd_ram_mem3_220_26, 
        p_wishbone_bd_ram_mem3_220_27, p_wishbone_bd_ram_mem3_220_28, 
        p_wishbone_bd_ram_mem3_220_29, p_wishbone_bd_ram_mem3_220_30, 
        p_wishbone_bd_ram_mem3_220_31, p_wishbone_bd_ram_mem3_221_24, 
        p_wishbone_bd_ram_mem3_221_25, p_wishbone_bd_ram_mem3_221_26, 
        p_wishbone_bd_ram_mem3_221_27, p_wishbone_bd_ram_mem3_221_28, 
        p_wishbone_bd_ram_mem3_221_29, p_wishbone_bd_ram_mem3_221_30, 
        p_wishbone_bd_ram_mem3_221_31, p_wishbone_bd_ram_mem3_222_24, 
        p_wishbone_bd_ram_mem3_222_25, p_wishbone_bd_ram_mem3_222_26, 
        p_wishbone_bd_ram_mem3_222_27, p_wishbone_bd_ram_mem3_222_28, 
        p_wishbone_bd_ram_mem3_222_29, p_wishbone_bd_ram_mem3_222_30, 
        p_wishbone_bd_ram_mem3_222_31, p_wishbone_bd_ram_mem3_223_24, 
        p_wishbone_bd_ram_mem3_223_25, p_wishbone_bd_ram_mem3_223_26, 
        p_wishbone_bd_ram_mem3_223_27, p_wishbone_bd_ram_mem3_223_28, 
        p_wishbone_bd_ram_mem3_223_29, p_wishbone_bd_ram_mem3_223_30, 
        p_wishbone_bd_ram_mem3_223_31, p_wishbone_bd_ram_mem3_224_24, 
        p_wishbone_bd_ram_mem3_224_25, p_wishbone_bd_ram_mem3_224_26, 
        p_wishbone_bd_ram_mem3_224_27, p_wishbone_bd_ram_mem3_224_28, 
        p_wishbone_bd_ram_mem3_224_29, p_wishbone_bd_ram_mem3_224_30, 
        p_wishbone_bd_ram_mem3_224_31, p_wishbone_bd_ram_mem3_225_24, 
        p_wishbone_bd_ram_mem3_225_25, p_wishbone_bd_ram_mem3_225_26, 
        p_wishbone_bd_ram_mem3_225_27, p_wishbone_bd_ram_mem3_225_28, 
        p_wishbone_bd_ram_mem3_225_29, p_wishbone_bd_ram_mem3_225_30, 
        p_wishbone_bd_ram_mem3_225_31, p_wishbone_bd_ram_mem3_226_24, 
        p_wishbone_bd_ram_mem3_226_25, p_wishbone_bd_ram_mem3_226_26, 
        p_wishbone_bd_ram_mem3_226_27, p_wishbone_bd_ram_mem3_226_28, 
        p_wishbone_bd_ram_mem3_226_29, p_wishbone_bd_ram_mem3_226_30, 
        p_wishbone_bd_ram_mem3_226_31, p_wishbone_bd_ram_mem3_227_24, 
        p_wishbone_bd_ram_mem3_227_25, p_wishbone_bd_ram_mem3_227_26, 
        p_wishbone_bd_ram_mem3_227_27, p_wishbone_bd_ram_mem3_227_28, 
        p_wishbone_bd_ram_mem3_227_29, p_wishbone_bd_ram_mem3_227_30, 
        p_wishbone_bd_ram_mem3_227_31, p_wishbone_bd_ram_mem3_228_24, 
        p_wishbone_bd_ram_mem3_228_25, p_wishbone_bd_ram_mem3_228_26, 
        p_wishbone_bd_ram_mem3_228_27, p_wishbone_bd_ram_mem3_228_28, 
        p_wishbone_bd_ram_mem3_228_29, p_wishbone_bd_ram_mem3_228_30, 
        p_wishbone_bd_ram_mem3_228_31, p_wishbone_bd_ram_mem3_229_24, 
        p_wishbone_bd_ram_mem3_229_25, p_wishbone_bd_ram_mem3_229_26, 
        p_wishbone_bd_ram_mem3_229_27, p_wishbone_bd_ram_mem3_229_28, 
        p_wishbone_bd_ram_mem3_229_29, p_wishbone_bd_ram_mem3_229_30, 
        p_wishbone_bd_ram_mem3_229_31, p_wishbone_bd_ram_mem3_230_24, 
        p_wishbone_bd_ram_mem3_230_25, p_wishbone_bd_ram_mem3_230_26, 
        p_wishbone_bd_ram_mem3_230_27, p_wishbone_bd_ram_mem3_230_28, 
        p_wishbone_bd_ram_mem3_230_29, p_wishbone_bd_ram_mem3_230_30, 
        p_wishbone_bd_ram_mem3_230_31, p_wishbone_bd_ram_mem3_231_24, 
        p_wishbone_bd_ram_mem3_231_25, p_wishbone_bd_ram_mem3_231_26, 
        p_wishbone_bd_ram_mem3_231_27, p_wishbone_bd_ram_mem3_231_28, 
        p_wishbone_bd_ram_mem3_231_29, p_wishbone_bd_ram_mem3_231_30, 
        p_wishbone_bd_ram_mem3_231_31, p_wishbone_bd_ram_mem3_232_24, 
        p_wishbone_bd_ram_mem3_232_25, p_wishbone_bd_ram_mem3_232_26, 
        p_wishbone_bd_ram_mem3_232_27, p_wishbone_bd_ram_mem3_232_28, 
        p_wishbone_bd_ram_mem3_232_29, p_wishbone_bd_ram_mem3_232_30, 
        p_wishbone_bd_ram_mem3_232_31, p_wishbone_bd_ram_mem3_233_24, 
        p_wishbone_bd_ram_mem3_233_25, p_wishbone_bd_ram_mem3_233_26, 
        p_wishbone_bd_ram_mem3_233_27, p_wishbone_bd_ram_mem3_233_28, 
        p_wishbone_bd_ram_mem3_233_29, p_wishbone_bd_ram_mem3_233_30, 
        p_wishbone_bd_ram_mem3_233_31, p_wishbone_bd_ram_mem3_234_24, 
        p_wishbone_bd_ram_mem3_234_25, p_wishbone_bd_ram_mem3_234_26, 
        p_wishbone_bd_ram_mem3_234_27, p_wishbone_bd_ram_mem3_234_28, 
        p_wishbone_bd_ram_mem3_234_29, p_wishbone_bd_ram_mem3_234_30, 
        p_wishbone_bd_ram_mem3_234_31, p_wishbone_bd_ram_mem3_235_24, 
        p_wishbone_bd_ram_mem3_235_25, p_wishbone_bd_ram_mem3_235_26, 
        p_wishbone_bd_ram_mem3_235_27, p_wishbone_bd_ram_mem3_235_28, 
        p_wishbone_bd_ram_mem3_235_29, p_wishbone_bd_ram_mem3_235_30, 
        p_wishbone_bd_ram_mem3_235_31, p_wishbone_bd_ram_mem3_236_24, 
        p_wishbone_bd_ram_mem3_236_25, p_wishbone_bd_ram_mem3_236_26, 
        p_wishbone_bd_ram_mem3_236_27, p_wishbone_bd_ram_mem3_236_28, 
        p_wishbone_bd_ram_mem3_236_29, p_wishbone_bd_ram_mem3_236_30, 
        p_wishbone_bd_ram_mem3_236_31, p_wishbone_bd_ram_mem3_237_24, 
        p_wishbone_bd_ram_mem3_237_25, p_wishbone_bd_ram_mem3_237_26, 
        p_wishbone_bd_ram_mem3_237_27, p_wishbone_bd_ram_mem3_237_28, 
        p_wishbone_bd_ram_mem3_237_29, p_wishbone_bd_ram_mem3_237_30, 
        p_wishbone_bd_ram_mem3_237_31, p_wishbone_bd_ram_mem3_238_24, 
        p_wishbone_bd_ram_mem3_238_25, p_wishbone_bd_ram_mem3_238_26, 
        p_wishbone_bd_ram_mem3_238_27, p_wishbone_bd_ram_mem3_238_28, 
        p_wishbone_bd_ram_mem3_238_29, p_wishbone_bd_ram_mem3_238_30, 
        p_wishbone_bd_ram_mem3_238_31, p_wishbone_bd_ram_mem3_239_24, 
        p_wishbone_bd_ram_mem3_239_25, p_wishbone_bd_ram_mem3_239_26, 
        p_wishbone_bd_ram_mem3_239_27, p_wishbone_bd_ram_mem3_239_28, 
        p_wishbone_bd_ram_mem3_239_29, p_wishbone_bd_ram_mem3_239_30, 
        p_wishbone_bd_ram_mem3_239_31, p_wishbone_bd_ram_mem3_240_24, 
        p_wishbone_bd_ram_mem3_240_25, p_wishbone_bd_ram_mem3_240_26, 
        p_wishbone_bd_ram_mem3_240_27, p_wishbone_bd_ram_mem3_240_28, 
        p_wishbone_bd_ram_mem3_240_29, p_wishbone_bd_ram_mem3_240_30, 
        p_wishbone_bd_ram_mem3_240_31, p_wishbone_bd_ram_mem3_241_24, 
        p_wishbone_bd_ram_mem3_241_25, p_wishbone_bd_ram_mem3_241_26, 
        p_wishbone_bd_ram_mem3_241_27, p_wishbone_bd_ram_mem3_241_28, 
        p_wishbone_bd_ram_mem3_241_29, p_wishbone_bd_ram_mem3_241_30, 
        p_wishbone_bd_ram_mem3_241_31, p_wishbone_bd_ram_mem3_242_24, 
        p_wishbone_bd_ram_mem3_242_25, p_wishbone_bd_ram_mem3_242_26, 
        p_wishbone_bd_ram_mem3_242_27, p_wishbone_bd_ram_mem3_242_28, 
        p_wishbone_bd_ram_mem3_242_29, p_wishbone_bd_ram_mem3_242_30, 
        p_wishbone_bd_ram_mem3_242_31, p_wishbone_bd_ram_mem3_243_24, 
        p_wishbone_bd_ram_mem3_243_25, p_wishbone_bd_ram_mem3_243_26, 
        p_wishbone_bd_ram_mem3_243_27, p_wishbone_bd_ram_mem3_243_28, 
        p_wishbone_bd_ram_mem3_243_29, p_wishbone_bd_ram_mem3_243_30, 
        p_wishbone_bd_ram_mem3_243_31, p_wishbone_bd_ram_mem3_244_24, 
        p_wishbone_bd_ram_mem3_244_25, p_wishbone_bd_ram_mem3_244_26, 
        p_wishbone_bd_ram_mem3_244_27, p_wishbone_bd_ram_mem3_244_28, 
        p_wishbone_bd_ram_mem3_244_29, p_wishbone_bd_ram_mem3_244_30, 
        p_wishbone_bd_ram_mem3_244_31, p_wishbone_bd_ram_mem3_245_24, 
        p_wishbone_bd_ram_mem3_245_25, p_wishbone_bd_ram_mem3_245_26, 
        p_wishbone_bd_ram_mem3_245_27, p_wishbone_bd_ram_mem3_245_28, 
        p_wishbone_bd_ram_mem3_245_29, p_wishbone_bd_ram_mem3_245_30, 
        p_wishbone_bd_ram_mem3_245_31, p_wishbone_bd_ram_mem3_246_24, 
        p_wishbone_bd_ram_mem3_246_25, p_wishbone_bd_ram_mem3_246_26, 
        p_wishbone_bd_ram_mem3_246_27, p_wishbone_bd_ram_mem3_246_28, 
        p_wishbone_bd_ram_mem3_246_29, p_wishbone_bd_ram_mem3_246_30, 
        p_wishbone_bd_ram_mem3_246_31, p_wishbone_bd_ram_mem3_247_24, 
        p_wishbone_bd_ram_mem3_247_25, p_wishbone_bd_ram_mem3_247_26, 
        p_wishbone_bd_ram_mem3_247_27, p_wishbone_bd_ram_mem3_247_28, 
        p_wishbone_bd_ram_mem3_247_29, p_wishbone_bd_ram_mem3_247_30, 
        p_wishbone_bd_ram_mem3_247_31, p_wishbone_bd_ram_mem3_248_24, 
        p_wishbone_bd_ram_mem3_248_25, p_wishbone_bd_ram_mem3_248_26, 
        p_wishbone_bd_ram_mem3_248_27, p_wishbone_bd_ram_mem3_248_28, 
        p_wishbone_bd_ram_mem3_248_29, p_wishbone_bd_ram_mem3_248_30, 
        p_wishbone_bd_ram_mem3_248_31, p_wishbone_bd_ram_mem3_249_24, 
        p_wishbone_bd_ram_mem3_249_25, p_wishbone_bd_ram_mem3_249_26, 
        p_wishbone_bd_ram_mem3_249_27, p_wishbone_bd_ram_mem3_249_28, 
        p_wishbone_bd_ram_mem3_249_29, p_wishbone_bd_ram_mem3_249_30, 
        p_wishbone_bd_ram_mem3_249_31, p_wishbone_bd_ram_mem3_250_24, 
        p_wishbone_bd_ram_mem3_250_25, p_wishbone_bd_ram_mem3_250_26, 
        p_wishbone_bd_ram_mem3_250_27, p_wishbone_bd_ram_mem3_250_28, 
        p_wishbone_bd_ram_mem3_250_29, p_wishbone_bd_ram_mem3_250_30, 
        p_wishbone_bd_ram_mem3_250_31, p_wishbone_bd_ram_mem3_251_24, 
        p_wishbone_bd_ram_mem3_251_25, p_wishbone_bd_ram_mem3_251_26, 
        p_wishbone_bd_ram_mem3_251_27, p_wishbone_bd_ram_mem3_251_28, 
        p_wishbone_bd_ram_mem3_251_29, p_wishbone_bd_ram_mem3_251_30, 
        p_wishbone_bd_ram_mem3_251_31, p_wishbone_bd_ram_mem3_252_24, 
        p_wishbone_bd_ram_mem3_252_25, p_wishbone_bd_ram_mem3_252_26, 
        p_wishbone_bd_ram_mem3_252_27, p_wishbone_bd_ram_mem3_252_28, 
        p_wishbone_bd_ram_mem3_252_29, p_wishbone_bd_ram_mem3_252_30, 
        p_wishbone_bd_ram_mem3_252_31, p_wishbone_bd_ram_mem3_253_24, 
        p_wishbone_bd_ram_mem3_253_25, p_wishbone_bd_ram_mem3_253_26, 
        p_wishbone_bd_ram_mem3_253_27, p_wishbone_bd_ram_mem3_253_28, 
        p_wishbone_bd_ram_mem3_253_29, p_wishbone_bd_ram_mem3_253_30, 
        p_wishbone_bd_ram_mem3_253_31, p_wishbone_bd_ram_mem3_254_24, 
        p_wishbone_bd_ram_mem3_254_25, p_wishbone_bd_ram_mem3_254_26, 
        p_wishbone_bd_ram_mem3_254_27, p_wishbone_bd_ram_mem3_254_28, 
        p_wishbone_bd_ram_mem3_254_29, p_wishbone_bd_ram_mem3_254_30, 
        p_wishbone_bd_ram_mem3_254_31, p_wishbone_bd_ram_mem3_255_24, 
        p_wishbone_bd_ram_mem3_255_25, p_wishbone_bd_ram_mem3_255_26, 
        p_wishbone_bd_ram_mem3_255_27, p_wishbone_bd_ram_mem3_255_28, 
        p_wishbone_bd_ram_mem3_255_29, p_wishbone_bd_ram_mem3_255_30, 
        p_wishbone_bd_ram_mem3_255_31, p_wishbone_bd_ram_mem1_0_8, 
        p_wishbone_bd_ram_mem1_0_9, p_wishbone_bd_ram_mem1_0_10, 
        p_wishbone_bd_ram_mem1_0_11, p_wishbone_bd_ram_mem1_0_12, 
        p_wishbone_bd_ram_mem1_0_13, p_wishbone_bd_ram_mem1_0_14, 
        p_wishbone_bd_ram_mem1_0_15, p_wishbone_bd_ram_mem1_1_8, 
        p_wishbone_bd_ram_mem1_1_9, p_wishbone_bd_ram_mem1_1_10, 
        p_wishbone_bd_ram_mem1_1_11, p_wishbone_bd_ram_mem1_1_12, 
        p_wishbone_bd_ram_mem1_1_13, p_wishbone_bd_ram_mem1_1_14, 
        p_wishbone_bd_ram_mem1_1_15, p_wishbone_bd_ram_mem1_2_8, 
        p_wishbone_bd_ram_mem1_2_9, p_wishbone_bd_ram_mem1_2_10, 
        p_wishbone_bd_ram_mem1_2_11, p_wishbone_bd_ram_mem1_2_12, 
        p_wishbone_bd_ram_mem1_2_13, p_wishbone_bd_ram_mem1_2_14, 
        p_wishbone_bd_ram_mem1_2_15, p_wishbone_bd_ram_mem1_3_8, 
        p_wishbone_bd_ram_mem1_3_9, p_wishbone_bd_ram_mem1_3_10, 
        p_wishbone_bd_ram_mem1_3_11, p_wishbone_bd_ram_mem1_3_12, 
        p_wishbone_bd_ram_mem1_3_13, p_wishbone_bd_ram_mem1_3_14, 
        p_wishbone_bd_ram_mem1_3_15, p_wishbone_bd_ram_mem1_4_8, 
        p_wishbone_bd_ram_mem1_4_9, p_wishbone_bd_ram_mem1_4_10, 
        p_wishbone_bd_ram_mem1_4_11, p_wishbone_bd_ram_mem1_4_12, 
        p_wishbone_bd_ram_mem1_4_13, p_wishbone_bd_ram_mem1_4_14, 
        p_wishbone_bd_ram_mem1_4_15, p_wishbone_bd_ram_mem1_5_8, 
        p_wishbone_bd_ram_mem1_5_9, p_wishbone_bd_ram_mem1_5_10, 
        p_wishbone_bd_ram_mem1_5_11, p_wishbone_bd_ram_mem1_5_12, 
        p_wishbone_bd_ram_mem1_5_13, p_wishbone_bd_ram_mem1_5_14, 
        p_wishbone_bd_ram_mem1_5_15, p_wishbone_bd_ram_mem1_6_8, 
        p_wishbone_bd_ram_mem1_6_9, p_wishbone_bd_ram_mem1_6_10, 
        p_wishbone_bd_ram_mem1_6_11, p_wishbone_bd_ram_mem1_6_12, 
        p_wishbone_bd_ram_mem1_6_13, p_wishbone_bd_ram_mem1_6_14, 
        p_wishbone_bd_ram_mem1_6_15, p_wishbone_bd_ram_mem1_7_8, 
        p_wishbone_bd_ram_mem1_7_9, p_wishbone_bd_ram_mem1_7_10, 
        p_wishbone_bd_ram_mem1_7_11, p_wishbone_bd_ram_mem1_7_12, 
        p_wishbone_bd_ram_mem1_7_13, p_wishbone_bd_ram_mem1_7_14, 
        p_wishbone_bd_ram_mem1_7_15, p_wishbone_bd_ram_mem1_8_8, 
        p_wishbone_bd_ram_mem1_8_9, p_wishbone_bd_ram_mem1_8_10, 
        p_wishbone_bd_ram_mem1_8_11, p_wishbone_bd_ram_mem1_8_12, 
        p_wishbone_bd_ram_mem1_8_13, p_wishbone_bd_ram_mem1_8_14, 
        p_wishbone_bd_ram_mem1_8_15, p_wishbone_bd_ram_mem1_9_8, 
        p_wishbone_bd_ram_mem1_9_9, p_wishbone_bd_ram_mem1_9_10, 
        p_wishbone_bd_ram_mem1_9_11, p_wishbone_bd_ram_mem1_9_12, 
        p_wishbone_bd_ram_mem1_9_13, p_wishbone_bd_ram_mem1_9_14, 
        p_wishbone_bd_ram_mem1_9_15, p_wishbone_bd_ram_mem1_10_8, 
        p_wishbone_bd_ram_mem1_10_9, p_wishbone_bd_ram_mem1_10_10, 
        p_wishbone_bd_ram_mem1_10_11, p_wishbone_bd_ram_mem1_10_12, 
        p_wishbone_bd_ram_mem1_10_13, p_wishbone_bd_ram_mem1_10_14, 
        p_wishbone_bd_ram_mem1_10_15, p_wishbone_bd_ram_mem1_11_8, 
        p_wishbone_bd_ram_mem1_11_9, p_wishbone_bd_ram_mem1_11_10, 
        p_wishbone_bd_ram_mem1_11_11, p_wishbone_bd_ram_mem1_11_12, 
        p_wishbone_bd_ram_mem1_11_13, p_wishbone_bd_ram_mem1_11_14, 
        p_wishbone_bd_ram_mem1_11_15, p_wishbone_bd_ram_mem1_12_8, 
        p_wishbone_bd_ram_mem1_12_9, p_wishbone_bd_ram_mem1_12_10, 
        p_wishbone_bd_ram_mem1_12_11, p_wishbone_bd_ram_mem1_12_12, 
        p_wishbone_bd_ram_mem1_12_13, p_wishbone_bd_ram_mem1_12_14, 
        p_wishbone_bd_ram_mem1_12_15, p_wishbone_bd_ram_mem1_13_8, 
        p_wishbone_bd_ram_mem1_13_9, p_wishbone_bd_ram_mem1_13_10, 
        p_wishbone_bd_ram_mem1_13_11, p_wishbone_bd_ram_mem1_13_12, 
        p_wishbone_bd_ram_mem1_13_13, p_wishbone_bd_ram_mem1_13_14, 
        p_wishbone_bd_ram_mem1_13_15, p_wishbone_bd_ram_mem1_14_8, 
        p_wishbone_bd_ram_mem1_14_9, p_wishbone_bd_ram_mem1_14_10, 
        p_wishbone_bd_ram_mem1_14_11, p_wishbone_bd_ram_mem1_14_12, 
        p_wishbone_bd_ram_mem1_14_13, p_wishbone_bd_ram_mem1_14_14, 
        p_wishbone_bd_ram_mem1_14_15, p_wishbone_bd_ram_mem1_15_8, 
        p_wishbone_bd_ram_mem1_15_9, p_wishbone_bd_ram_mem1_15_10, 
        p_wishbone_bd_ram_mem1_15_11, p_wishbone_bd_ram_mem1_15_12, 
        p_wishbone_bd_ram_mem1_15_13, p_wishbone_bd_ram_mem1_15_14, 
        p_wishbone_bd_ram_mem1_15_15, p_wishbone_bd_ram_mem1_16_8, 
        p_wishbone_bd_ram_mem1_16_9, p_wishbone_bd_ram_mem1_16_10, 
        p_wishbone_bd_ram_mem1_16_11, p_wishbone_bd_ram_mem1_16_12, 
        p_wishbone_bd_ram_mem1_16_13, p_wishbone_bd_ram_mem1_16_14, 
        p_wishbone_bd_ram_mem1_16_15, p_wishbone_bd_ram_mem1_17_8, 
        p_wishbone_bd_ram_mem1_17_9, p_wishbone_bd_ram_mem1_17_10, 
        p_wishbone_bd_ram_mem1_17_11, p_wishbone_bd_ram_mem1_17_12, 
        p_wishbone_bd_ram_mem1_17_13, p_wishbone_bd_ram_mem1_17_14, 
        p_wishbone_bd_ram_mem1_17_15, p_wishbone_bd_ram_mem1_18_8, 
        p_wishbone_bd_ram_mem1_18_9, p_wishbone_bd_ram_mem1_18_10, 
        p_wishbone_bd_ram_mem1_18_11, p_wishbone_bd_ram_mem1_18_12, 
        p_wishbone_bd_ram_mem1_18_13, p_wishbone_bd_ram_mem1_18_14, 
        p_wishbone_bd_ram_mem1_18_15, p_wishbone_bd_ram_mem1_19_8, 
        p_wishbone_bd_ram_mem1_19_9, p_wishbone_bd_ram_mem1_19_10, 
        p_wishbone_bd_ram_mem1_19_11, p_wishbone_bd_ram_mem1_19_12, 
        p_wishbone_bd_ram_mem1_19_13, p_wishbone_bd_ram_mem1_19_14, 
        p_wishbone_bd_ram_mem1_19_15, p_wishbone_bd_ram_mem1_20_8, 
        p_wishbone_bd_ram_mem1_20_9, p_wishbone_bd_ram_mem1_20_10, 
        p_wishbone_bd_ram_mem1_20_11, p_wishbone_bd_ram_mem1_20_12, 
        p_wishbone_bd_ram_mem1_20_13, p_wishbone_bd_ram_mem1_20_14, 
        p_wishbone_bd_ram_mem1_20_15, p_wishbone_bd_ram_mem1_21_8, 
        p_wishbone_bd_ram_mem1_21_9, p_wishbone_bd_ram_mem1_21_10, 
        p_wishbone_bd_ram_mem1_21_11, p_wishbone_bd_ram_mem1_21_12, 
        p_wishbone_bd_ram_mem1_21_13, p_wishbone_bd_ram_mem1_21_14, 
        p_wishbone_bd_ram_mem1_21_15, p_wishbone_bd_ram_mem1_22_8, 
        p_wishbone_bd_ram_mem1_22_9, p_wishbone_bd_ram_mem1_22_10, 
        p_wishbone_bd_ram_mem1_22_11, p_wishbone_bd_ram_mem1_22_12, 
        p_wishbone_bd_ram_mem1_22_13, p_wishbone_bd_ram_mem1_22_14, 
        p_wishbone_bd_ram_mem1_22_15, p_wishbone_bd_ram_mem1_23_8, 
        p_wishbone_bd_ram_mem1_23_9, p_wishbone_bd_ram_mem1_23_10, 
        p_wishbone_bd_ram_mem1_23_11, p_wishbone_bd_ram_mem1_23_12, 
        p_wishbone_bd_ram_mem1_23_13, p_wishbone_bd_ram_mem1_23_14, 
        p_wishbone_bd_ram_mem1_23_15, p_wishbone_bd_ram_mem1_24_8, 
        p_wishbone_bd_ram_mem1_24_9, p_wishbone_bd_ram_mem1_24_10, 
        p_wishbone_bd_ram_mem1_24_11, p_wishbone_bd_ram_mem1_24_12, 
        p_wishbone_bd_ram_mem1_24_13, p_wishbone_bd_ram_mem1_24_14, 
        p_wishbone_bd_ram_mem1_24_15, p_wishbone_bd_ram_mem1_25_8, 
        p_wishbone_bd_ram_mem1_25_9, p_wishbone_bd_ram_mem1_25_10, 
        p_wishbone_bd_ram_mem1_25_11, p_wishbone_bd_ram_mem1_25_12, 
        p_wishbone_bd_ram_mem1_25_13, p_wishbone_bd_ram_mem1_25_14, 
        p_wishbone_bd_ram_mem1_25_15, p_wishbone_bd_ram_mem1_26_8, 
        p_wishbone_bd_ram_mem1_26_9, p_wishbone_bd_ram_mem1_26_10, 
        p_wishbone_bd_ram_mem1_26_11, p_wishbone_bd_ram_mem1_26_12, 
        p_wishbone_bd_ram_mem1_26_13, p_wishbone_bd_ram_mem1_26_14, 
        p_wishbone_bd_ram_mem1_26_15, p_wishbone_bd_ram_mem1_27_8, 
        p_wishbone_bd_ram_mem1_27_9, p_wishbone_bd_ram_mem1_27_10, 
        p_wishbone_bd_ram_mem1_27_11, p_wishbone_bd_ram_mem1_27_12, 
        p_wishbone_bd_ram_mem1_27_13, p_wishbone_bd_ram_mem1_27_14, 
        p_wishbone_bd_ram_mem1_27_15, p_wishbone_bd_ram_mem1_28_8, 
        p_wishbone_bd_ram_mem1_28_9, p_wishbone_bd_ram_mem1_28_10, 
        p_wishbone_bd_ram_mem1_28_11, p_wishbone_bd_ram_mem1_28_12, 
        p_wishbone_bd_ram_mem1_28_13, p_wishbone_bd_ram_mem1_28_14, 
        p_wishbone_bd_ram_mem1_28_15, p_wishbone_bd_ram_mem1_29_8, 
        p_wishbone_bd_ram_mem1_29_9, p_wishbone_bd_ram_mem1_29_10, 
        p_wishbone_bd_ram_mem1_29_11, p_wishbone_bd_ram_mem1_29_12, 
        p_wishbone_bd_ram_mem1_29_13, p_wishbone_bd_ram_mem1_29_14, 
        p_wishbone_bd_ram_mem1_29_15, p_wishbone_bd_ram_mem1_30_8, 
        p_wishbone_bd_ram_mem1_30_9, p_wishbone_bd_ram_mem1_30_10, 
        p_wishbone_bd_ram_mem1_30_11, p_wishbone_bd_ram_mem1_30_12, 
        p_wishbone_bd_ram_mem1_30_13, p_wishbone_bd_ram_mem1_30_14, 
        p_wishbone_bd_ram_mem1_30_15, p_wishbone_bd_ram_mem1_31_8, 
        p_wishbone_bd_ram_mem1_31_9, p_wishbone_bd_ram_mem1_31_10, 
        p_wishbone_bd_ram_mem1_31_11, p_wishbone_bd_ram_mem1_31_12, 
        p_wishbone_bd_ram_mem1_31_13, p_wishbone_bd_ram_mem1_31_14, 
        p_wishbone_bd_ram_mem1_31_15, p_wishbone_bd_ram_mem1_32_8, 
        p_wishbone_bd_ram_mem1_32_9, p_wishbone_bd_ram_mem1_32_10, 
        p_wishbone_bd_ram_mem1_32_11, p_wishbone_bd_ram_mem1_32_12, 
        p_wishbone_bd_ram_mem1_32_13, p_wishbone_bd_ram_mem1_32_14, 
        p_wishbone_bd_ram_mem1_32_15, p_wishbone_bd_ram_mem1_33_8, 
        p_wishbone_bd_ram_mem1_33_9, p_wishbone_bd_ram_mem1_33_10, 
        p_wishbone_bd_ram_mem1_33_11, p_wishbone_bd_ram_mem1_33_12, 
        p_wishbone_bd_ram_mem1_33_13, p_wishbone_bd_ram_mem1_33_14, 
        p_wishbone_bd_ram_mem1_33_15, p_wishbone_bd_ram_mem1_34_8, 
        p_wishbone_bd_ram_mem1_34_9, p_wishbone_bd_ram_mem1_34_10, 
        p_wishbone_bd_ram_mem1_34_11, p_wishbone_bd_ram_mem1_34_12, 
        p_wishbone_bd_ram_mem1_34_13, p_wishbone_bd_ram_mem1_34_14, 
        p_wishbone_bd_ram_mem1_34_15, p_wishbone_bd_ram_mem1_35_8, 
        p_wishbone_bd_ram_mem1_35_9, p_wishbone_bd_ram_mem1_35_10, 
        p_wishbone_bd_ram_mem1_35_11, p_wishbone_bd_ram_mem1_35_12, 
        p_wishbone_bd_ram_mem1_35_13, p_wishbone_bd_ram_mem1_35_14, 
        p_wishbone_bd_ram_mem1_35_15, p_wishbone_bd_ram_mem1_36_8, 
        p_wishbone_bd_ram_mem1_36_9, p_wishbone_bd_ram_mem1_36_10, 
        p_wishbone_bd_ram_mem1_36_11, p_wishbone_bd_ram_mem1_36_12, 
        p_wishbone_bd_ram_mem1_36_13, p_wishbone_bd_ram_mem1_36_14, 
        p_wishbone_bd_ram_mem1_36_15, p_wishbone_bd_ram_mem1_37_8, 
        p_wishbone_bd_ram_mem1_37_9, p_wishbone_bd_ram_mem1_37_10, 
        p_wishbone_bd_ram_mem1_37_11, p_wishbone_bd_ram_mem1_37_12, 
        p_wishbone_bd_ram_mem1_37_13, p_wishbone_bd_ram_mem1_37_14, 
        p_wishbone_bd_ram_mem1_37_15, p_wishbone_bd_ram_mem1_38_8, 
        p_wishbone_bd_ram_mem1_38_9, p_wishbone_bd_ram_mem1_38_10, 
        p_wishbone_bd_ram_mem1_38_11, p_wishbone_bd_ram_mem1_38_12, 
        p_wishbone_bd_ram_mem1_38_13, p_wishbone_bd_ram_mem1_38_14, 
        p_wishbone_bd_ram_mem1_38_15, p_wishbone_bd_ram_mem1_39_8, 
        p_wishbone_bd_ram_mem1_39_9, p_wishbone_bd_ram_mem1_39_10, 
        p_wishbone_bd_ram_mem1_39_11, p_wishbone_bd_ram_mem1_39_12, 
        p_wishbone_bd_ram_mem1_39_13, p_wishbone_bd_ram_mem1_39_14, 
        p_wishbone_bd_ram_mem1_39_15, p_wishbone_bd_ram_mem1_40_8, 
        p_wishbone_bd_ram_mem1_40_9, p_wishbone_bd_ram_mem1_40_10, 
        p_wishbone_bd_ram_mem1_40_11, p_wishbone_bd_ram_mem1_40_12, 
        p_wishbone_bd_ram_mem1_40_13, p_wishbone_bd_ram_mem1_40_14, 
        p_wishbone_bd_ram_mem1_40_15, p_wishbone_bd_ram_mem1_41_8, 
        p_wishbone_bd_ram_mem1_41_9, p_wishbone_bd_ram_mem1_41_10, 
        p_wishbone_bd_ram_mem1_41_11, p_wishbone_bd_ram_mem1_41_12, 
        p_wishbone_bd_ram_mem1_41_13, p_wishbone_bd_ram_mem1_41_14, 
        p_wishbone_bd_ram_mem1_41_15, p_wishbone_bd_ram_mem1_42_8, 
        p_wishbone_bd_ram_mem1_42_9, p_wishbone_bd_ram_mem1_42_10, 
        p_wishbone_bd_ram_mem1_42_11, p_wishbone_bd_ram_mem1_42_12, 
        p_wishbone_bd_ram_mem1_42_13, p_wishbone_bd_ram_mem1_42_14, 
        p_wishbone_bd_ram_mem1_42_15, p_wishbone_bd_ram_mem1_43_8, 
        p_wishbone_bd_ram_mem1_43_9, p_wishbone_bd_ram_mem1_43_10, 
        p_wishbone_bd_ram_mem1_43_11, p_wishbone_bd_ram_mem1_43_12, 
        p_wishbone_bd_ram_mem1_43_13, p_wishbone_bd_ram_mem1_43_14, 
        p_wishbone_bd_ram_mem1_43_15, p_wishbone_bd_ram_mem1_44_8, 
        p_wishbone_bd_ram_mem1_44_9, p_wishbone_bd_ram_mem1_44_10, 
        p_wishbone_bd_ram_mem1_44_11, p_wishbone_bd_ram_mem1_44_12, 
        p_wishbone_bd_ram_mem1_44_13, p_wishbone_bd_ram_mem1_44_14, 
        p_wishbone_bd_ram_mem1_44_15, p_wishbone_bd_ram_mem1_45_8, 
        p_wishbone_bd_ram_mem1_45_9, p_wishbone_bd_ram_mem1_45_10, 
        p_wishbone_bd_ram_mem1_45_11, p_wishbone_bd_ram_mem1_45_12, 
        p_wishbone_bd_ram_mem1_45_13, p_wishbone_bd_ram_mem1_45_14, 
        p_wishbone_bd_ram_mem1_45_15, p_wishbone_bd_ram_mem1_46_8, 
        p_wishbone_bd_ram_mem1_46_9, p_wishbone_bd_ram_mem1_46_10, 
        p_wishbone_bd_ram_mem1_46_11, p_wishbone_bd_ram_mem1_46_12, 
        p_wishbone_bd_ram_mem1_46_13, p_wishbone_bd_ram_mem1_46_14, 
        p_wishbone_bd_ram_mem1_46_15, p_wishbone_bd_ram_mem1_47_8, 
        p_wishbone_bd_ram_mem1_47_9, p_wishbone_bd_ram_mem1_47_10, 
        p_wishbone_bd_ram_mem1_47_11, p_wishbone_bd_ram_mem1_47_12, 
        p_wishbone_bd_ram_mem1_47_13, p_wishbone_bd_ram_mem1_47_14, 
        p_wishbone_bd_ram_mem1_47_15, p_wishbone_bd_ram_mem1_48_8, 
        p_wishbone_bd_ram_mem1_48_9, p_wishbone_bd_ram_mem1_48_10, 
        p_wishbone_bd_ram_mem1_48_11, p_wishbone_bd_ram_mem1_48_12, 
        p_wishbone_bd_ram_mem1_48_13, p_wishbone_bd_ram_mem1_48_14, 
        p_wishbone_bd_ram_mem1_48_15, p_wishbone_bd_ram_mem1_49_8, 
        p_wishbone_bd_ram_mem1_49_9, p_wishbone_bd_ram_mem1_49_10, 
        p_wishbone_bd_ram_mem1_49_11, p_wishbone_bd_ram_mem1_49_12, 
        p_wishbone_bd_ram_mem1_49_13, p_wishbone_bd_ram_mem1_49_14, 
        p_wishbone_bd_ram_mem1_49_15, p_wishbone_bd_ram_mem1_50_8, 
        p_wishbone_bd_ram_mem1_50_9, p_wishbone_bd_ram_mem1_50_10, 
        p_wishbone_bd_ram_mem1_50_11, p_wishbone_bd_ram_mem1_50_12, 
        p_wishbone_bd_ram_mem1_50_13, p_wishbone_bd_ram_mem1_50_14, 
        p_wishbone_bd_ram_mem1_50_15, p_wishbone_bd_ram_mem1_51_8, 
        p_wishbone_bd_ram_mem1_51_9, p_wishbone_bd_ram_mem1_51_10, 
        p_wishbone_bd_ram_mem1_51_11, p_wishbone_bd_ram_mem1_51_12, 
        p_wishbone_bd_ram_mem1_51_13, p_wishbone_bd_ram_mem1_51_14, 
        p_wishbone_bd_ram_mem1_51_15, p_wishbone_bd_ram_mem1_52_8, 
        p_wishbone_bd_ram_mem1_52_9, p_wishbone_bd_ram_mem1_52_10, 
        p_wishbone_bd_ram_mem1_52_11, p_wishbone_bd_ram_mem1_52_12, 
        p_wishbone_bd_ram_mem1_52_13, p_wishbone_bd_ram_mem1_52_14, 
        p_wishbone_bd_ram_mem1_52_15, p_wishbone_bd_ram_mem1_53_8, 
        p_wishbone_bd_ram_mem1_53_9, p_wishbone_bd_ram_mem1_53_10, 
        p_wishbone_bd_ram_mem1_53_11, p_wishbone_bd_ram_mem1_53_12, 
        p_wishbone_bd_ram_mem1_53_13, p_wishbone_bd_ram_mem1_53_14, 
        p_wishbone_bd_ram_mem1_53_15, p_wishbone_bd_ram_mem1_54_8, 
        p_wishbone_bd_ram_mem1_54_9, p_wishbone_bd_ram_mem1_54_10, 
        p_wishbone_bd_ram_mem1_54_11, p_wishbone_bd_ram_mem1_54_12, 
        p_wishbone_bd_ram_mem1_54_13, p_wishbone_bd_ram_mem1_54_14, 
        p_wishbone_bd_ram_mem1_54_15, p_wishbone_bd_ram_mem1_55_8, 
        p_wishbone_bd_ram_mem1_55_9, p_wishbone_bd_ram_mem1_55_10, 
        p_wishbone_bd_ram_mem1_55_11, p_wishbone_bd_ram_mem1_55_12, 
        p_wishbone_bd_ram_mem1_55_13, p_wishbone_bd_ram_mem1_55_14, 
        p_wishbone_bd_ram_mem1_55_15, p_wishbone_bd_ram_mem1_56_8, 
        p_wishbone_bd_ram_mem1_56_9, p_wishbone_bd_ram_mem1_56_10, 
        p_wishbone_bd_ram_mem1_56_11, p_wishbone_bd_ram_mem1_56_12, 
        p_wishbone_bd_ram_mem1_56_13, p_wishbone_bd_ram_mem1_56_14, 
        p_wishbone_bd_ram_mem1_56_15, p_wishbone_bd_ram_mem1_57_8, 
        p_wishbone_bd_ram_mem1_57_9, p_wishbone_bd_ram_mem1_57_10, 
        p_wishbone_bd_ram_mem1_57_11, p_wishbone_bd_ram_mem1_57_12, 
        p_wishbone_bd_ram_mem1_57_13, p_wishbone_bd_ram_mem1_57_14, 
        p_wishbone_bd_ram_mem1_57_15, p_wishbone_bd_ram_mem1_58_8, 
        p_wishbone_bd_ram_mem1_58_9, p_wishbone_bd_ram_mem1_58_10, 
        p_wishbone_bd_ram_mem1_58_11, p_wishbone_bd_ram_mem1_58_12, 
        p_wishbone_bd_ram_mem1_58_13, p_wishbone_bd_ram_mem1_58_14, 
        p_wishbone_bd_ram_mem1_58_15, p_wishbone_bd_ram_mem1_59_8, 
        p_wishbone_bd_ram_mem1_59_9, p_wishbone_bd_ram_mem1_59_10, 
        p_wishbone_bd_ram_mem1_59_11, p_wishbone_bd_ram_mem1_59_12, 
        p_wishbone_bd_ram_mem1_59_13, p_wishbone_bd_ram_mem1_59_14, 
        p_wishbone_bd_ram_mem1_59_15, p_wishbone_bd_ram_mem1_60_8, 
        p_wishbone_bd_ram_mem1_60_9, p_wishbone_bd_ram_mem1_60_10, 
        p_wishbone_bd_ram_mem1_60_11, p_wishbone_bd_ram_mem1_60_12, 
        p_wishbone_bd_ram_mem1_60_13, p_wishbone_bd_ram_mem1_60_14, 
        p_wishbone_bd_ram_mem1_60_15, p_wishbone_bd_ram_mem1_61_8, 
        p_wishbone_bd_ram_mem1_61_9, p_wishbone_bd_ram_mem1_61_10, 
        p_wishbone_bd_ram_mem1_61_11, p_wishbone_bd_ram_mem1_61_12, 
        p_wishbone_bd_ram_mem1_61_13, p_wishbone_bd_ram_mem1_61_14, 
        p_wishbone_bd_ram_mem1_61_15, p_wishbone_bd_ram_mem1_62_8, 
        p_wishbone_bd_ram_mem1_62_9, p_wishbone_bd_ram_mem1_62_10, 
        p_wishbone_bd_ram_mem1_62_11, p_wishbone_bd_ram_mem1_62_12, 
        p_wishbone_bd_ram_mem1_62_13, p_wishbone_bd_ram_mem1_62_14, 
        p_wishbone_bd_ram_mem1_62_15, p_wishbone_bd_ram_mem1_63_8, 
        p_wishbone_bd_ram_mem1_63_9, p_wishbone_bd_ram_mem1_63_10, 
        p_wishbone_bd_ram_mem1_63_11, p_wishbone_bd_ram_mem1_63_12, 
        p_wishbone_bd_ram_mem1_63_13, p_wishbone_bd_ram_mem1_63_14, 
        p_wishbone_bd_ram_mem1_63_15, p_wishbone_bd_ram_mem1_64_8, 
        p_wishbone_bd_ram_mem1_64_9, p_wishbone_bd_ram_mem1_64_10, 
        p_wishbone_bd_ram_mem1_64_11, p_wishbone_bd_ram_mem1_64_12, 
        p_wishbone_bd_ram_mem1_64_13, p_wishbone_bd_ram_mem1_64_14, 
        p_wishbone_bd_ram_mem1_64_15, p_wishbone_bd_ram_mem1_65_8, 
        p_wishbone_bd_ram_mem1_65_9, p_wishbone_bd_ram_mem1_65_10, 
        p_wishbone_bd_ram_mem1_65_11, p_wishbone_bd_ram_mem1_65_12, 
        p_wishbone_bd_ram_mem1_65_13, p_wishbone_bd_ram_mem1_65_14, 
        p_wishbone_bd_ram_mem1_65_15, p_wishbone_bd_ram_mem1_66_8, 
        p_wishbone_bd_ram_mem1_66_9, p_wishbone_bd_ram_mem1_66_10, 
        p_wishbone_bd_ram_mem1_66_11, p_wishbone_bd_ram_mem1_66_12, 
        p_wishbone_bd_ram_mem1_66_13, p_wishbone_bd_ram_mem1_66_14, 
        p_wishbone_bd_ram_mem1_66_15, p_wishbone_bd_ram_mem1_67_8, 
        p_wishbone_bd_ram_mem1_67_9, p_wishbone_bd_ram_mem1_67_10, 
        p_wishbone_bd_ram_mem1_67_11, p_wishbone_bd_ram_mem1_67_12, 
        p_wishbone_bd_ram_mem1_67_13, p_wishbone_bd_ram_mem1_67_14, 
        p_wishbone_bd_ram_mem1_67_15, p_wishbone_bd_ram_mem1_68_8, 
        p_wishbone_bd_ram_mem1_68_9, p_wishbone_bd_ram_mem1_68_10, 
        p_wishbone_bd_ram_mem1_68_11, p_wishbone_bd_ram_mem1_68_12, 
        p_wishbone_bd_ram_mem1_68_13, p_wishbone_bd_ram_mem1_68_14, 
        p_wishbone_bd_ram_mem1_68_15, p_wishbone_bd_ram_mem1_69_8, 
        p_wishbone_bd_ram_mem1_69_9, p_wishbone_bd_ram_mem1_69_10, 
        p_wishbone_bd_ram_mem1_69_11, p_wishbone_bd_ram_mem1_69_12, 
        p_wishbone_bd_ram_mem1_69_13, p_wishbone_bd_ram_mem1_69_14, 
        p_wishbone_bd_ram_mem1_69_15, p_wishbone_bd_ram_mem1_70_8, 
        p_wishbone_bd_ram_mem1_70_9, p_wishbone_bd_ram_mem1_70_10, 
        p_wishbone_bd_ram_mem1_70_11, p_wishbone_bd_ram_mem1_70_12, 
        p_wishbone_bd_ram_mem1_70_13, p_wishbone_bd_ram_mem1_70_14, 
        p_wishbone_bd_ram_mem1_70_15, p_wishbone_bd_ram_mem1_71_8, 
        p_wishbone_bd_ram_mem1_71_9, p_wishbone_bd_ram_mem1_71_10, 
        p_wishbone_bd_ram_mem1_71_11, p_wishbone_bd_ram_mem1_71_12, 
        p_wishbone_bd_ram_mem1_71_13, p_wishbone_bd_ram_mem1_71_14, 
        p_wishbone_bd_ram_mem1_71_15, p_wishbone_bd_ram_mem1_72_8, 
        p_wishbone_bd_ram_mem1_72_9, p_wishbone_bd_ram_mem1_72_10, 
        p_wishbone_bd_ram_mem1_72_11, p_wishbone_bd_ram_mem1_72_12, 
        p_wishbone_bd_ram_mem1_72_13, p_wishbone_bd_ram_mem1_72_14, 
        p_wishbone_bd_ram_mem1_72_15, p_wishbone_bd_ram_mem1_73_8, 
        p_wishbone_bd_ram_mem1_73_9, p_wishbone_bd_ram_mem1_73_10, 
        p_wishbone_bd_ram_mem1_73_11, p_wishbone_bd_ram_mem1_73_12, 
        p_wishbone_bd_ram_mem1_73_13, p_wishbone_bd_ram_mem1_73_14, 
        p_wishbone_bd_ram_mem1_73_15, p_wishbone_bd_ram_mem1_74_8, 
        p_wishbone_bd_ram_mem1_74_9, p_wishbone_bd_ram_mem1_74_10, 
        p_wishbone_bd_ram_mem1_74_11, p_wishbone_bd_ram_mem1_74_12, 
        p_wishbone_bd_ram_mem1_74_13, p_wishbone_bd_ram_mem1_74_14, 
        p_wishbone_bd_ram_mem1_74_15, p_wishbone_bd_ram_mem1_75_8, 
        p_wishbone_bd_ram_mem1_75_9, p_wishbone_bd_ram_mem1_75_10, 
        p_wishbone_bd_ram_mem1_75_11, p_wishbone_bd_ram_mem1_75_12, 
        p_wishbone_bd_ram_mem1_75_13, p_wishbone_bd_ram_mem1_75_14, 
        p_wishbone_bd_ram_mem1_75_15, p_wishbone_bd_ram_mem1_76_8, 
        p_wishbone_bd_ram_mem1_76_9, p_wishbone_bd_ram_mem1_76_10, 
        p_wishbone_bd_ram_mem1_76_11, p_wishbone_bd_ram_mem1_76_12, 
        p_wishbone_bd_ram_mem1_76_13, p_wishbone_bd_ram_mem1_76_14, 
        p_wishbone_bd_ram_mem1_76_15, p_wishbone_bd_ram_mem1_77_8, 
        p_wishbone_bd_ram_mem1_77_9, p_wishbone_bd_ram_mem1_77_10, 
        p_wishbone_bd_ram_mem1_77_11, p_wishbone_bd_ram_mem1_77_12, 
        p_wishbone_bd_ram_mem1_77_13, p_wishbone_bd_ram_mem1_77_14, 
        p_wishbone_bd_ram_mem1_77_15, p_wishbone_bd_ram_mem1_78_8, 
        p_wishbone_bd_ram_mem1_78_9, p_wishbone_bd_ram_mem1_78_10, 
        p_wishbone_bd_ram_mem1_78_11, p_wishbone_bd_ram_mem1_78_12, 
        p_wishbone_bd_ram_mem1_78_13, p_wishbone_bd_ram_mem1_78_14, 
        p_wishbone_bd_ram_mem1_78_15, p_wishbone_bd_ram_mem1_79_8, 
        p_wishbone_bd_ram_mem1_79_9, p_wishbone_bd_ram_mem1_79_10, 
        p_wishbone_bd_ram_mem1_79_11, p_wishbone_bd_ram_mem1_79_12, 
        p_wishbone_bd_ram_mem1_79_13, p_wishbone_bd_ram_mem1_79_14, 
        p_wishbone_bd_ram_mem1_79_15, p_wishbone_bd_ram_mem1_80_8, 
        p_wishbone_bd_ram_mem1_80_9, p_wishbone_bd_ram_mem1_80_10, 
        p_wishbone_bd_ram_mem1_80_11, p_wishbone_bd_ram_mem1_80_12, 
        p_wishbone_bd_ram_mem1_80_13, p_wishbone_bd_ram_mem1_80_14, 
        p_wishbone_bd_ram_mem1_80_15, p_wishbone_bd_ram_mem1_81_8, 
        p_wishbone_bd_ram_mem1_81_9, p_wishbone_bd_ram_mem1_81_10, 
        p_wishbone_bd_ram_mem1_81_11, p_wishbone_bd_ram_mem1_81_12, 
        p_wishbone_bd_ram_mem1_81_13, p_wishbone_bd_ram_mem1_81_14, 
        p_wishbone_bd_ram_mem1_81_15, p_wishbone_bd_ram_mem1_82_8, 
        p_wishbone_bd_ram_mem1_82_9, p_wishbone_bd_ram_mem1_82_10, 
        p_wishbone_bd_ram_mem1_82_11, p_wishbone_bd_ram_mem1_82_12, 
        p_wishbone_bd_ram_mem1_82_13, p_wishbone_bd_ram_mem1_82_14, 
        p_wishbone_bd_ram_mem1_82_15, p_wishbone_bd_ram_mem1_83_8, 
        p_wishbone_bd_ram_mem1_83_9, p_wishbone_bd_ram_mem1_83_10, 
        p_wishbone_bd_ram_mem1_83_11, p_wishbone_bd_ram_mem1_83_12, 
        p_wishbone_bd_ram_mem1_83_13, p_wishbone_bd_ram_mem1_83_14, 
        p_wishbone_bd_ram_mem1_83_15, p_wishbone_bd_ram_mem1_84_8, 
        p_wishbone_bd_ram_mem1_84_9, p_wishbone_bd_ram_mem1_84_10, 
        p_wishbone_bd_ram_mem1_84_11, p_wishbone_bd_ram_mem1_84_12, 
        p_wishbone_bd_ram_mem1_84_13, p_wishbone_bd_ram_mem1_84_14, 
        p_wishbone_bd_ram_mem1_84_15, p_wishbone_bd_ram_mem1_85_8, 
        p_wishbone_bd_ram_mem1_85_9, p_wishbone_bd_ram_mem1_85_10, 
        p_wishbone_bd_ram_mem1_85_11, p_wishbone_bd_ram_mem1_85_12, 
        p_wishbone_bd_ram_mem1_85_13, p_wishbone_bd_ram_mem1_85_14, 
        p_wishbone_bd_ram_mem1_85_15, p_wishbone_bd_ram_mem1_86_8, 
        p_wishbone_bd_ram_mem1_86_9, p_wishbone_bd_ram_mem1_86_10, 
        p_wishbone_bd_ram_mem1_86_11, p_wishbone_bd_ram_mem1_86_12, 
        p_wishbone_bd_ram_mem1_86_13, p_wishbone_bd_ram_mem1_86_14, 
        p_wishbone_bd_ram_mem1_86_15, p_wishbone_bd_ram_mem1_87_8, 
        p_wishbone_bd_ram_mem1_87_9, p_wishbone_bd_ram_mem1_87_10, 
        p_wishbone_bd_ram_mem1_87_11, p_wishbone_bd_ram_mem1_87_12, 
        p_wishbone_bd_ram_mem1_87_13, p_wishbone_bd_ram_mem1_87_14, 
        p_wishbone_bd_ram_mem1_87_15, p_wishbone_bd_ram_mem1_88_8, 
        p_wishbone_bd_ram_mem1_88_9, p_wishbone_bd_ram_mem1_88_10, 
        p_wishbone_bd_ram_mem1_88_11, p_wishbone_bd_ram_mem1_88_12, 
        p_wishbone_bd_ram_mem1_88_13, p_wishbone_bd_ram_mem1_88_14, 
        p_wishbone_bd_ram_mem1_88_15, p_wishbone_bd_ram_mem1_89_8, 
        p_wishbone_bd_ram_mem1_89_9, p_wishbone_bd_ram_mem1_89_10, 
        p_wishbone_bd_ram_mem1_89_11, p_wishbone_bd_ram_mem1_89_12, 
        p_wishbone_bd_ram_mem1_89_13, p_wishbone_bd_ram_mem1_89_14, 
        p_wishbone_bd_ram_mem1_89_15, p_wishbone_bd_ram_mem1_90_8, 
        p_wishbone_bd_ram_mem1_90_9, p_wishbone_bd_ram_mem1_90_10, 
        p_wishbone_bd_ram_mem1_90_11, p_wishbone_bd_ram_mem1_90_12, 
        p_wishbone_bd_ram_mem1_90_13, p_wishbone_bd_ram_mem1_90_14, 
        p_wishbone_bd_ram_mem1_90_15, p_wishbone_bd_ram_mem1_91_8, 
        p_wishbone_bd_ram_mem1_91_9, p_wishbone_bd_ram_mem1_91_10, 
        p_wishbone_bd_ram_mem1_91_11, p_wishbone_bd_ram_mem1_91_12, 
        p_wishbone_bd_ram_mem1_91_13, p_wishbone_bd_ram_mem1_91_14, 
        p_wishbone_bd_ram_mem1_91_15, p_wishbone_bd_ram_mem1_92_8, 
        p_wishbone_bd_ram_mem1_92_9, p_wishbone_bd_ram_mem1_92_10, 
        p_wishbone_bd_ram_mem1_92_11, p_wishbone_bd_ram_mem1_92_12, 
        p_wishbone_bd_ram_mem1_92_13, p_wishbone_bd_ram_mem1_92_14, 
        p_wishbone_bd_ram_mem1_92_15, p_wishbone_bd_ram_mem1_93_8, 
        p_wishbone_bd_ram_mem1_93_9, p_wishbone_bd_ram_mem1_93_10, 
        p_wishbone_bd_ram_mem1_93_11, p_wishbone_bd_ram_mem1_93_12, 
        p_wishbone_bd_ram_mem1_93_13, p_wishbone_bd_ram_mem1_93_14, 
        p_wishbone_bd_ram_mem1_93_15, p_wishbone_bd_ram_mem1_94_8, 
        p_wishbone_bd_ram_mem1_94_9, p_wishbone_bd_ram_mem1_94_10, 
        p_wishbone_bd_ram_mem1_94_11, p_wishbone_bd_ram_mem1_94_12, 
        p_wishbone_bd_ram_mem1_94_13, p_wishbone_bd_ram_mem1_94_14, 
        p_wishbone_bd_ram_mem1_94_15, p_wishbone_bd_ram_mem1_95_8, 
        p_wishbone_bd_ram_mem1_95_9, p_wishbone_bd_ram_mem1_95_10, 
        p_wishbone_bd_ram_mem1_95_11, p_wishbone_bd_ram_mem1_95_12, 
        p_wishbone_bd_ram_mem1_95_13, p_wishbone_bd_ram_mem1_95_14, 
        p_wishbone_bd_ram_mem1_95_15, p_wishbone_bd_ram_mem1_96_8, 
        p_wishbone_bd_ram_mem1_96_9, p_wishbone_bd_ram_mem1_96_10, 
        p_wishbone_bd_ram_mem1_96_11, p_wishbone_bd_ram_mem1_96_12, 
        p_wishbone_bd_ram_mem1_96_13, p_wishbone_bd_ram_mem1_96_14, 
        p_wishbone_bd_ram_mem1_96_15, p_wishbone_bd_ram_mem1_97_8, 
        p_wishbone_bd_ram_mem1_97_9, p_wishbone_bd_ram_mem1_97_10, 
        p_wishbone_bd_ram_mem1_97_11, p_wishbone_bd_ram_mem1_97_12, 
        p_wishbone_bd_ram_mem1_97_13, p_wishbone_bd_ram_mem1_97_14, 
        p_wishbone_bd_ram_mem1_97_15, p_wishbone_bd_ram_mem1_98_8, 
        p_wishbone_bd_ram_mem1_98_9, p_wishbone_bd_ram_mem1_98_10, 
        p_wishbone_bd_ram_mem1_98_11, p_wishbone_bd_ram_mem1_98_12, 
        p_wishbone_bd_ram_mem1_98_13, p_wishbone_bd_ram_mem1_98_14, 
        p_wishbone_bd_ram_mem1_98_15, p_wishbone_bd_ram_mem1_99_8, 
        p_wishbone_bd_ram_mem1_99_9, p_wishbone_bd_ram_mem1_99_10, 
        p_wishbone_bd_ram_mem1_99_11, p_wishbone_bd_ram_mem1_99_12, 
        p_wishbone_bd_ram_mem1_99_13, p_wishbone_bd_ram_mem1_99_14, 
        p_wishbone_bd_ram_mem1_99_15, p_wishbone_bd_ram_mem1_100_8, 
        p_wishbone_bd_ram_mem1_100_9, p_wishbone_bd_ram_mem1_100_10, 
        p_wishbone_bd_ram_mem1_100_11, p_wishbone_bd_ram_mem1_100_12, 
        p_wishbone_bd_ram_mem1_100_13, p_wishbone_bd_ram_mem1_100_14, 
        p_wishbone_bd_ram_mem1_100_15, p_wishbone_bd_ram_mem1_101_8, 
        p_wishbone_bd_ram_mem1_101_9, p_wishbone_bd_ram_mem1_101_10, 
        p_wishbone_bd_ram_mem1_101_11, p_wishbone_bd_ram_mem1_101_12, 
        p_wishbone_bd_ram_mem1_101_13, p_wishbone_bd_ram_mem1_101_14, 
        p_wishbone_bd_ram_mem1_101_15, p_wishbone_bd_ram_mem1_102_8, 
        p_wishbone_bd_ram_mem1_102_9, p_wishbone_bd_ram_mem1_102_10, 
        p_wishbone_bd_ram_mem1_102_11, p_wishbone_bd_ram_mem1_102_12, 
        p_wishbone_bd_ram_mem1_102_13, p_wishbone_bd_ram_mem1_102_14, 
        p_wishbone_bd_ram_mem1_102_15, p_wishbone_bd_ram_mem1_103_8, 
        p_wishbone_bd_ram_mem1_103_9, p_wishbone_bd_ram_mem1_103_10, 
        p_wishbone_bd_ram_mem1_103_11, p_wishbone_bd_ram_mem1_103_12, 
        p_wishbone_bd_ram_mem1_103_13, p_wishbone_bd_ram_mem1_103_14, 
        p_wishbone_bd_ram_mem1_103_15, p_wishbone_bd_ram_mem1_104_8, 
        p_wishbone_bd_ram_mem1_104_9, p_wishbone_bd_ram_mem1_104_10, 
        p_wishbone_bd_ram_mem1_104_11, p_wishbone_bd_ram_mem1_104_12, 
        p_wishbone_bd_ram_mem1_104_13, p_wishbone_bd_ram_mem1_104_14, 
        p_wishbone_bd_ram_mem1_104_15, p_wishbone_bd_ram_mem1_105_8, 
        p_wishbone_bd_ram_mem1_105_9, p_wishbone_bd_ram_mem1_105_10, 
        p_wishbone_bd_ram_mem1_105_11, p_wishbone_bd_ram_mem1_105_12, 
        p_wishbone_bd_ram_mem1_105_13, p_wishbone_bd_ram_mem1_105_14, 
        p_wishbone_bd_ram_mem1_105_15, p_wishbone_bd_ram_mem1_106_8, 
        p_wishbone_bd_ram_mem1_106_9, p_wishbone_bd_ram_mem1_106_10, 
        p_wishbone_bd_ram_mem1_106_11, p_wishbone_bd_ram_mem1_106_12, 
        p_wishbone_bd_ram_mem1_106_13, p_wishbone_bd_ram_mem1_106_14, 
        p_wishbone_bd_ram_mem1_106_15, p_wishbone_bd_ram_mem1_107_8, 
        p_wishbone_bd_ram_mem1_107_9, p_wishbone_bd_ram_mem1_107_10, 
        p_wishbone_bd_ram_mem1_107_11, p_wishbone_bd_ram_mem1_107_12, 
        p_wishbone_bd_ram_mem1_107_13, p_wishbone_bd_ram_mem1_107_14, 
        p_wishbone_bd_ram_mem1_107_15, p_wishbone_bd_ram_mem1_108_8, 
        p_wishbone_bd_ram_mem1_108_9, p_wishbone_bd_ram_mem1_108_10, 
        p_wishbone_bd_ram_mem1_108_11, p_wishbone_bd_ram_mem1_108_12, 
        p_wishbone_bd_ram_mem1_108_13, p_wishbone_bd_ram_mem1_108_14, 
        p_wishbone_bd_ram_mem1_108_15, p_wishbone_bd_ram_mem1_109_8, 
        p_wishbone_bd_ram_mem1_109_9, p_wishbone_bd_ram_mem1_109_10, 
        p_wishbone_bd_ram_mem1_109_11, p_wishbone_bd_ram_mem1_109_12, 
        p_wishbone_bd_ram_mem1_109_13, p_wishbone_bd_ram_mem1_109_14, 
        p_wishbone_bd_ram_mem1_109_15, p_wishbone_bd_ram_mem1_110_8, 
        p_wishbone_bd_ram_mem1_110_9, p_wishbone_bd_ram_mem1_110_10, 
        p_wishbone_bd_ram_mem1_110_11, p_wishbone_bd_ram_mem1_110_12, 
        p_wishbone_bd_ram_mem1_110_13, p_wishbone_bd_ram_mem1_110_14, 
        p_wishbone_bd_ram_mem1_110_15, p_wishbone_bd_ram_mem1_111_8, 
        p_wishbone_bd_ram_mem1_111_9, p_wishbone_bd_ram_mem1_111_10, 
        p_wishbone_bd_ram_mem1_111_11, p_wishbone_bd_ram_mem1_111_12, 
        p_wishbone_bd_ram_mem1_111_13, p_wishbone_bd_ram_mem1_111_14, 
        p_wishbone_bd_ram_mem1_111_15, p_wishbone_bd_ram_mem1_112_8, 
        p_wishbone_bd_ram_mem1_112_9, p_wishbone_bd_ram_mem1_112_10, 
        p_wishbone_bd_ram_mem1_112_11, p_wishbone_bd_ram_mem1_112_12, 
        p_wishbone_bd_ram_mem1_112_13, p_wishbone_bd_ram_mem1_112_14, 
        p_wishbone_bd_ram_mem1_112_15, p_wishbone_bd_ram_mem1_113_8, 
        p_wishbone_bd_ram_mem1_113_9, p_wishbone_bd_ram_mem1_113_10, 
        p_wishbone_bd_ram_mem1_113_11, p_wishbone_bd_ram_mem1_113_12, 
        p_wishbone_bd_ram_mem1_113_13, p_wishbone_bd_ram_mem1_113_14, 
        p_wishbone_bd_ram_mem1_113_15, p_wishbone_bd_ram_mem1_114_8, 
        p_wishbone_bd_ram_mem1_114_9, p_wishbone_bd_ram_mem1_114_10, 
        p_wishbone_bd_ram_mem1_114_11, p_wishbone_bd_ram_mem1_114_12, 
        p_wishbone_bd_ram_mem1_114_13, p_wishbone_bd_ram_mem1_114_14, 
        p_wishbone_bd_ram_mem1_114_15, p_wishbone_bd_ram_mem1_115_8, 
        p_wishbone_bd_ram_mem1_115_9, p_wishbone_bd_ram_mem1_115_10, 
        p_wishbone_bd_ram_mem1_115_11, p_wishbone_bd_ram_mem1_115_12, 
        p_wishbone_bd_ram_mem1_115_13, p_wishbone_bd_ram_mem1_115_14, 
        p_wishbone_bd_ram_mem1_115_15, p_wishbone_bd_ram_mem1_116_8, 
        p_wishbone_bd_ram_mem1_116_9, p_wishbone_bd_ram_mem1_116_10, 
        p_wishbone_bd_ram_mem1_116_11, p_wishbone_bd_ram_mem1_116_12, 
        p_wishbone_bd_ram_mem1_116_13, p_wishbone_bd_ram_mem1_116_14, 
        p_wishbone_bd_ram_mem1_116_15, p_wishbone_bd_ram_mem1_117_8, 
        p_wishbone_bd_ram_mem1_117_9, p_wishbone_bd_ram_mem1_117_10, 
        p_wishbone_bd_ram_mem1_117_11, p_wishbone_bd_ram_mem1_117_12, 
        p_wishbone_bd_ram_mem1_117_13, p_wishbone_bd_ram_mem1_117_14, 
        p_wishbone_bd_ram_mem1_117_15, p_wishbone_bd_ram_mem1_118_8, 
        p_wishbone_bd_ram_mem1_118_9, p_wishbone_bd_ram_mem1_118_10, 
        p_wishbone_bd_ram_mem1_118_11, p_wishbone_bd_ram_mem1_118_12, 
        p_wishbone_bd_ram_mem1_118_13, p_wishbone_bd_ram_mem1_118_14, 
        p_wishbone_bd_ram_mem1_118_15, p_wishbone_bd_ram_mem1_119_8, 
        p_wishbone_bd_ram_mem1_119_9, p_wishbone_bd_ram_mem1_119_10, 
        p_wishbone_bd_ram_mem1_119_11, p_wishbone_bd_ram_mem1_119_12, 
        p_wishbone_bd_ram_mem1_119_13, p_wishbone_bd_ram_mem1_119_14, 
        p_wishbone_bd_ram_mem1_119_15, p_wishbone_bd_ram_mem1_120_8, 
        p_wishbone_bd_ram_mem1_120_9, p_wishbone_bd_ram_mem1_120_10, 
        p_wishbone_bd_ram_mem1_120_11, p_wishbone_bd_ram_mem1_120_12, 
        p_wishbone_bd_ram_mem1_120_13, p_wishbone_bd_ram_mem1_120_14, 
        p_wishbone_bd_ram_mem1_120_15, p_wishbone_bd_ram_mem1_121_8, 
        p_wishbone_bd_ram_mem1_121_9, p_wishbone_bd_ram_mem1_121_10, 
        p_wishbone_bd_ram_mem1_121_11, p_wishbone_bd_ram_mem1_121_12, 
        p_wishbone_bd_ram_mem1_121_13, p_wishbone_bd_ram_mem1_121_14, 
        p_wishbone_bd_ram_mem1_121_15, p_wishbone_bd_ram_mem1_122_8, 
        p_wishbone_bd_ram_mem1_122_9, p_wishbone_bd_ram_mem1_122_10, 
        p_wishbone_bd_ram_mem1_122_11, p_wishbone_bd_ram_mem1_122_12, 
        p_wishbone_bd_ram_mem1_122_13, p_wishbone_bd_ram_mem1_122_14, 
        p_wishbone_bd_ram_mem1_122_15, p_wishbone_bd_ram_mem1_123_8, 
        p_wishbone_bd_ram_mem1_123_9, p_wishbone_bd_ram_mem1_123_10, 
        p_wishbone_bd_ram_mem1_123_11, p_wishbone_bd_ram_mem1_123_12, 
        p_wishbone_bd_ram_mem1_123_13, p_wishbone_bd_ram_mem1_123_14, 
        p_wishbone_bd_ram_mem1_123_15, p_wishbone_bd_ram_mem1_124_8, 
        p_wishbone_bd_ram_mem1_124_9, p_wishbone_bd_ram_mem1_124_10, 
        p_wishbone_bd_ram_mem1_124_11, p_wishbone_bd_ram_mem1_124_12, 
        p_wishbone_bd_ram_mem1_124_13, p_wishbone_bd_ram_mem1_124_14, 
        p_wishbone_bd_ram_mem1_124_15, p_wishbone_bd_ram_mem1_125_8, 
        p_wishbone_bd_ram_mem1_125_9, p_wishbone_bd_ram_mem1_125_10, 
        p_wishbone_bd_ram_mem1_125_11, p_wishbone_bd_ram_mem1_125_12, 
        p_wishbone_bd_ram_mem1_125_13, p_wishbone_bd_ram_mem1_125_14, 
        p_wishbone_bd_ram_mem1_125_15, p_wishbone_bd_ram_mem1_126_8, 
        p_wishbone_bd_ram_mem1_126_9, p_wishbone_bd_ram_mem1_126_10, 
        p_wishbone_bd_ram_mem1_126_11, p_wishbone_bd_ram_mem1_126_12, 
        p_wishbone_bd_ram_mem1_126_13, p_wishbone_bd_ram_mem1_126_14, 
        p_wishbone_bd_ram_mem1_126_15, p_wishbone_bd_ram_mem1_127_8, 
        p_wishbone_bd_ram_mem1_127_9, p_wishbone_bd_ram_mem1_127_10, 
        p_wishbone_bd_ram_mem1_127_11, p_wishbone_bd_ram_mem1_127_12, 
        p_wishbone_bd_ram_mem1_127_13, p_wishbone_bd_ram_mem1_127_14, 
        p_wishbone_bd_ram_mem1_127_15, p_wishbone_bd_ram_mem1_128_8, 
        p_wishbone_bd_ram_mem1_128_9, p_wishbone_bd_ram_mem1_128_10, 
        p_wishbone_bd_ram_mem1_128_11, p_wishbone_bd_ram_mem1_128_12, 
        p_wishbone_bd_ram_mem1_128_13, p_wishbone_bd_ram_mem1_128_14, 
        p_wishbone_bd_ram_mem1_128_15, p_wishbone_bd_ram_mem1_129_8, 
        p_wishbone_bd_ram_mem1_129_9, p_wishbone_bd_ram_mem1_129_10, 
        p_wishbone_bd_ram_mem1_129_11, p_wishbone_bd_ram_mem1_129_12, 
        p_wishbone_bd_ram_mem1_129_13, p_wishbone_bd_ram_mem1_129_14, 
        p_wishbone_bd_ram_mem1_129_15, p_wishbone_bd_ram_mem1_130_8, 
        p_wishbone_bd_ram_mem1_130_9, p_wishbone_bd_ram_mem1_130_10, 
        p_wishbone_bd_ram_mem1_130_11, p_wishbone_bd_ram_mem1_130_12, 
        p_wishbone_bd_ram_mem1_130_13, p_wishbone_bd_ram_mem1_130_14, 
        p_wishbone_bd_ram_mem1_130_15, p_wishbone_bd_ram_mem1_131_8, 
        p_wishbone_bd_ram_mem1_131_9, p_wishbone_bd_ram_mem1_131_10, 
        p_wishbone_bd_ram_mem1_131_11, p_wishbone_bd_ram_mem1_131_12, 
        p_wishbone_bd_ram_mem1_131_13, p_wishbone_bd_ram_mem1_131_14, 
        p_wishbone_bd_ram_mem1_131_15, p_wishbone_bd_ram_mem1_132_8, 
        p_wishbone_bd_ram_mem1_132_9, p_wishbone_bd_ram_mem1_132_10, 
        p_wishbone_bd_ram_mem1_132_11, p_wishbone_bd_ram_mem1_132_12, 
        p_wishbone_bd_ram_mem1_132_13, p_wishbone_bd_ram_mem1_132_14, 
        p_wishbone_bd_ram_mem1_132_15, p_wishbone_bd_ram_mem1_133_8, 
        p_wishbone_bd_ram_mem1_133_9, p_wishbone_bd_ram_mem1_133_10, 
        p_wishbone_bd_ram_mem1_133_11, p_wishbone_bd_ram_mem1_133_12, 
        p_wishbone_bd_ram_mem1_133_13, p_wishbone_bd_ram_mem1_133_14, 
        p_wishbone_bd_ram_mem1_133_15, p_wishbone_bd_ram_mem1_134_8, 
        p_wishbone_bd_ram_mem1_134_9, p_wishbone_bd_ram_mem1_134_10, 
        p_wishbone_bd_ram_mem1_134_11, p_wishbone_bd_ram_mem1_134_12, 
        p_wishbone_bd_ram_mem1_134_13, p_wishbone_bd_ram_mem1_134_14, 
        p_wishbone_bd_ram_mem1_134_15, p_wishbone_bd_ram_mem1_135_8, 
        p_wishbone_bd_ram_mem1_135_9, p_wishbone_bd_ram_mem1_135_10, 
        p_wishbone_bd_ram_mem1_135_11, p_wishbone_bd_ram_mem1_135_12, 
        p_wishbone_bd_ram_mem1_135_13, p_wishbone_bd_ram_mem1_135_14, 
        p_wishbone_bd_ram_mem1_135_15, p_wishbone_bd_ram_mem1_136_8, 
        p_wishbone_bd_ram_mem1_136_9, p_wishbone_bd_ram_mem1_136_10, 
        p_wishbone_bd_ram_mem1_136_11, p_wishbone_bd_ram_mem1_136_12, 
        p_wishbone_bd_ram_mem1_136_13, p_wishbone_bd_ram_mem1_136_14, 
        p_wishbone_bd_ram_mem1_136_15, p_wishbone_bd_ram_mem1_137_8, 
        p_wishbone_bd_ram_mem1_137_9, p_wishbone_bd_ram_mem1_137_10, 
        p_wishbone_bd_ram_mem1_137_11, p_wishbone_bd_ram_mem1_137_12, 
        p_wishbone_bd_ram_mem1_137_13, p_wishbone_bd_ram_mem1_137_14, 
        p_wishbone_bd_ram_mem1_137_15, p_wishbone_bd_ram_mem1_138_8, 
        p_wishbone_bd_ram_mem1_138_9, p_wishbone_bd_ram_mem1_138_10, 
        p_wishbone_bd_ram_mem1_138_11, p_wishbone_bd_ram_mem1_138_12, 
        p_wishbone_bd_ram_mem1_138_13, p_wishbone_bd_ram_mem1_138_14, 
        p_wishbone_bd_ram_mem1_138_15, p_wishbone_bd_ram_mem1_139_8, 
        p_wishbone_bd_ram_mem1_139_9, p_wishbone_bd_ram_mem1_139_10, 
        p_wishbone_bd_ram_mem1_139_11, p_wishbone_bd_ram_mem1_139_12, 
        p_wishbone_bd_ram_mem1_139_13, p_wishbone_bd_ram_mem1_139_14, 
        p_wishbone_bd_ram_mem1_139_15, p_wishbone_bd_ram_mem1_140_8, 
        p_wishbone_bd_ram_mem1_140_9, p_wishbone_bd_ram_mem1_140_10, 
        p_wishbone_bd_ram_mem1_140_11, p_wishbone_bd_ram_mem1_140_12, 
        p_wishbone_bd_ram_mem1_140_13, p_wishbone_bd_ram_mem1_140_14, 
        p_wishbone_bd_ram_mem1_140_15, p_wishbone_bd_ram_mem1_141_8, 
        p_wishbone_bd_ram_mem1_141_9, p_wishbone_bd_ram_mem1_141_10, 
        p_wishbone_bd_ram_mem1_141_11, p_wishbone_bd_ram_mem1_141_12, 
        p_wishbone_bd_ram_mem1_141_13, p_wishbone_bd_ram_mem1_141_14, 
        p_wishbone_bd_ram_mem1_141_15, p_wishbone_bd_ram_mem1_142_8, 
        p_wishbone_bd_ram_mem1_142_9, p_wishbone_bd_ram_mem1_142_10, 
        p_wishbone_bd_ram_mem1_142_11, p_wishbone_bd_ram_mem1_142_12, 
        p_wishbone_bd_ram_mem1_142_13, p_wishbone_bd_ram_mem1_142_14, 
        p_wishbone_bd_ram_mem1_142_15, p_wishbone_bd_ram_mem1_143_8, 
        p_wishbone_bd_ram_mem1_143_9, p_wishbone_bd_ram_mem1_143_10, 
        p_wishbone_bd_ram_mem1_143_11, p_wishbone_bd_ram_mem1_143_12, 
        p_wishbone_bd_ram_mem1_143_13, p_wishbone_bd_ram_mem1_143_14, 
        p_wishbone_bd_ram_mem1_143_15, p_wishbone_bd_ram_mem1_144_8, 
        p_wishbone_bd_ram_mem1_144_9, p_wishbone_bd_ram_mem1_144_10, 
        p_wishbone_bd_ram_mem1_144_11, p_wishbone_bd_ram_mem1_144_12, 
        p_wishbone_bd_ram_mem1_144_13, p_wishbone_bd_ram_mem1_144_14, 
        p_wishbone_bd_ram_mem1_144_15, p_wishbone_bd_ram_mem1_145_8, 
        p_wishbone_bd_ram_mem1_145_9, p_wishbone_bd_ram_mem1_145_10, 
        p_wishbone_bd_ram_mem1_145_11, p_wishbone_bd_ram_mem1_145_12, 
        p_wishbone_bd_ram_mem1_145_13, p_wishbone_bd_ram_mem1_145_14, 
        p_wishbone_bd_ram_mem1_145_15, p_wishbone_bd_ram_mem1_146_8, 
        p_wishbone_bd_ram_mem1_146_9, p_wishbone_bd_ram_mem1_146_10, 
        p_wishbone_bd_ram_mem1_146_11, p_wishbone_bd_ram_mem1_146_12, 
        p_wishbone_bd_ram_mem1_146_13, p_wishbone_bd_ram_mem1_146_14, 
        p_wishbone_bd_ram_mem1_146_15, p_wishbone_bd_ram_mem1_147_8, 
        p_wishbone_bd_ram_mem1_147_9, p_wishbone_bd_ram_mem1_147_10, 
        p_wishbone_bd_ram_mem1_147_11, p_wishbone_bd_ram_mem1_147_12, 
        p_wishbone_bd_ram_mem1_147_13, p_wishbone_bd_ram_mem1_147_14, 
        p_wishbone_bd_ram_mem1_147_15, p_wishbone_bd_ram_mem1_148_8, 
        p_wishbone_bd_ram_mem1_148_9, p_wishbone_bd_ram_mem1_148_10, 
        p_wishbone_bd_ram_mem1_148_11, p_wishbone_bd_ram_mem1_148_12, 
        p_wishbone_bd_ram_mem1_148_13, p_wishbone_bd_ram_mem1_148_14, 
        p_wishbone_bd_ram_mem1_148_15, p_wishbone_bd_ram_mem1_149_8, 
        p_wishbone_bd_ram_mem1_149_9, p_wishbone_bd_ram_mem1_149_10, 
        p_wishbone_bd_ram_mem1_149_11, p_wishbone_bd_ram_mem1_149_12, 
        p_wishbone_bd_ram_mem1_149_13, p_wishbone_bd_ram_mem1_149_14, 
        p_wishbone_bd_ram_mem1_149_15, p_wishbone_bd_ram_mem1_150_8, 
        p_wishbone_bd_ram_mem1_150_9, p_wishbone_bd_ram_mem1_150_10, 
        p_wishbone_bd_ram_mem1_150_11, p_wishbone_bd_ram_mem1_150_12, 
        p_wishbone_bd_ram_mem1_150_13, p_wishbone_bd_ram_mem1_150_14, 
        p_wishbone_bd_ram_mem1_150_15, p_wishbone_bd_ram_mem1_151_8, 
        p_wishbone_bd_ram_mem1_151_9, p_wishbone_bd_ram_mem1_151_10, 
        p_wishbone_bd_ram_mem1_151_11, p_wishbone_bd_ram_mem1_151_12, 
        p_wishbone_bd_ram_mem1_151_13, p_wishbone_bd_ram_mem1_151_14, 
        p_wishbone_bd_ram_mem1_151_15, p_wishbone_bd_ram_mem1_152_8, 
        p_wishbone_bd_ram_mem1_152_9, p_wishbone_bd_ram_mem1_152_10, 
        p_wishbone_bd_ram_mem1_152_11, p_wishbone_bd_ram_mem1_152_12, 
        p_wishbone_bd_ram_mem1_152_13, p_wishbone_bd_ram_mem1_152_14, 
        p_wishbone_bd_ram_mem1_152_15, p_wishbone_bd_ram_mem1_153_8, 
        p_wishbone_bd_ram_mem1_153_9, p_wishbone_bd_ram_mem1_153_10, 
        p_wishbone_bd_ram_mem1_153_11, p_wishbone_bd_ram_mem1_153_12, 
        p_wishbone_bd_ram_mem1_153_13, p_wishbone_bd_ram_mem1_153_14, 
        p_wishbone_bd_ram_mem1_153_15, p_wishbone_bd_ram_mem1_154_8, 
        p_wishbone_bd_ram_mem1_154_9, p_wishbone_bd_ram_mem1_154_10, 
        p_wishbone_bd_ram_mem1_154_11, p_wishbone_bd_ram_mem1_154_12, 
        p_wishbone_bd_ram_mem1_154_13, p_wishbone_bd_ram_mem1_154_14, 
        p_wishbone_bd_ram_mem1_154_15, p_wishbone_bd_ram_mem1_155_8, 
        p_wishbone_bd_ram_mem1_155_9, p_wishbone_bd_ram_mem1_155_10, 
        p_wishbone_bd_ram_mem1_155_11, p_wishbone_bd_ram_mem1_155_12, 
        p_wishbone_bd_ram_mem1_155_13, p_wishbone_bd_ram_mem1_155_14, 
        p_wishbone_bd_ram_mem1_155_15, p_wishbone_bd_ram_mem1_156_8, 
        p_wishbone_bd_ram_mem1_156_9, p_wishbone_bd_ram_mem1_156_10, 
        p_wishbone_bd_ram_mem1_156_11, p_wishbone_bd_ram_mem1_156_12, 
        p_wishbone_bd_ram_mem1_156_13, p_wishbone_bd_ram_mem1_156_14, 
        p_wishbone_bd_ram_mem1_156_15, p_wishbone_bd_ram_mem1_157_8, 
        p_wishbone_bd_ram_mem1_157_9, p_wishbone_bd_ram_mem1_157_10, 
        p_wishbone_bd_ram_mem1_157_11, p_wishbone_bd_ram_mem1_157_12, 
        p_wishbone_bd_ram_mem1_157_13, p_wishbone_bd_ram_mem1_157_14, 
        p_wishbone_bd_ram_mem1_157_15, p_wishbone_bd_ram_mem1_158_8, 
        p_wishbone_bd_ram_mem1_158_9, p_wishbone_bd_ram_mem1_158_10, 
        p_wishbone_bd_ram_mem1_158_11, p_wishbone_bd_ram_mem1_158_12, 
        p_wishbone_bd_ram_mem1_158_13, p_wishbone_bd_ram_mem1_158_14, 
        p_wishbone_bd_ram_mem1_158_15, p_wishbone_bd_ram_mem1_159_8, 
        p_wishbone_bd_ram_mem1_159_9, p_wishbone_bd_ram_mem1_159_10, 
        p_wishbone_bd_ram_mem1_159_11, p_wishbone_bd_ram_mem1_159_12, 
        p_wishbone_bd_ram_mem1_159_13, p_wishbone_bd_ram_mem1_159_14, 
        p_wishbone_bd_ram_mem1_159_15, p_wishbone_bd_ram_mem1_160_8, 
        p_wishbone_bd_ram_mem1_160_9, p_wishbone_bd_ram_mem1_160_10, 
        p_wishbone_bd_ram_mem1_160_11, p_wishbone_bd_ram_mem1_160_12, 
        p_wishbone_bd_ram_mem1_160_13, p_wishbone_bd_ram_mem1_160_14, 
        p_wishbone_bd_ram_mem1_160_15, p_wishbone_bd_ram_mem1_161_8, 
        p_wishbone_bd_ram_mem1_161_9, p_wishbone_bd_ram_mem1_161_10, 
        p_wishbone_bd_ram_mem1_161_11, p_wishbone_bd_ram_mem1_161_12, 
        p_wishbone_bd_ram_mem1_161_13, p_wishbone_bd_ram_mem1_161_14, 
        p_wishbone_bd_ram_mem1_161_15, p_wishbone_bd_ram_mem1_162_8, 
        p_wishbone_bd_ram_mem1_162_9, p_wishbone_bd_ram_mem1_162_10, 
        p_wishbone_bd_ram_mem1_162_11, p_wishbone_bd_ram_mem1_162_12, 
        p_wishbone_bd_ram_mem1_162_13, p_wishbone_bd_ram_mem1_162_14, 
        p_wishbone_bd_ram_mem1_162_15, p_wishbone_bd_ram_mem1_163_8, 
        p_wishbone_bd_ram_mem1_163_9, p_wishbone_bd_ram_mem1_163_10, 
        p_wishbone_bd_ram_mem1_163_11, p_wishbone_bd_ram_mem1_163_12, 
        p_wishbone_bd_ram_mem1_163_13, p_wishbone_bd_ram_mem1_163_14, 
        p_wishbone_bd_ram_mem1_163_15, p_wishbone_bd_ram_mem1_164_8, 
        p_wishbone_bd_ram_mem1_164_9, p_wishbone_bd_ram_mem1_164_10, 
        p_wishbone_bd_ram_mem1_164_11, p_wishbone_bd_ram_mem1_164_12, 
        p_wishbone_bd_ram_mem1_164_13, p_wishbone_bd_ram_mem1_164_14, 
        p_wishbone_bd_ram_mem1_164_15, p_wishbone_bd_ram_mem1_165_8, 
        p_wishbone_bd_ram_mem1_165_9, p_wishbone_bd_ram_mem1_165_10, 
        p_wishbone_bd_ram_mem1_165_11, p_wishbone_bd_ram_mem1_165_12, 
        p_wishbone_bd_ram_mem1_165_13, p_wishbone_bd_ram_mem1_165_14, 
        p_wishbone_bd_ram_mem1_165_15, p_wishbone_bd_ram_mem1_166_8, 
        p_wishbone_bd_ram_mem1_166_9, p_wishbone_bd_ram_mem1_166_10, 
        p_wishbone_bd_ram_mem1_166_11, p_wishbone_bd_ram_mem1_166_12, 
        p_wishbone_bd_ram_mem1_166_13, p_wishbone_bd_ram_mem1_166_14, 
        p_wishbone_bd_ram_mem1_166_15, p_wishbone_bd_ram_mem1_167_8, 
        p_wishbone_bd_ram_mem1_167_9, p_wishbone_bd_ram_mem1_167_10, 
        p_wishbone_bd_ram_mem1_167_11, p_wishbone_bd_ram_mem1_167_12, 
        p_wishbone_bd_ram_mem1_167_13, p_wishbone_bd_ram_mem1_167_14, 
        p_wishbone_bd_ram_mem1_167_15, p_wishbone_bd_ram_mem1_168_8, 
        p_wishbone_bd_ram_mem1_168_9, p_wishbone_bd_ram_mem1_168_10, 
        p_wishbone_bd_ram_mem1_168_11, p_wishbone_bd_ram_mem1_168_12, 
        p_wishbone_bd_ram_mem1_168_13, p_wishbone_bd_ram_mem1_168_14, 
        p_wishbone_bd_ram_mem1_168_15, p_wishbone_bd_ram_mem1_169_8, 
        p_wishbone_bd_ram_mem1_169_9, p_wishbone_bd_ram_mem1_169_10, 
        p_wishbone_bd_ram_mem1_169_11, p_wishbone_bd_ram_mem1_169_12, 
        p_wishbone_bd_ram_mem1_169_13, p_wishbone_bd_ram_mem1_169_14, 
        p_wishbone_bd_ram_mem1_169_15, p_wishbone_bd_ram_mem1_170_8, 
        p_wishbone_bd_ram_mem1_170_9, p_wishbone_bd_ram_mem1_170_10, 
        p_wishbone_bd_ram_mem1_170_11, p_wishbone_bd_ram_mem1_170_12, 
        p_wishbone_bd_ram_mem1_170_13, p_wishbone_bd_ram_mem1_170_14, 
        p_wishbone_bd_ram_mem1_170_15, p_wishbone_bd_ram_mem1_171_8, 
        p_wishbone_bd_ram_mem1_171_9, p_wishbone_bd_ram_mem1_171_10, 
        p_wishbone_bd_ram_mem1_171_11, p_wishbone_bd_ram_mem1_171_12, 
        p_wishbone_bd_ram_mem1_171_13, p_wishbone_bd_ram_mem1_171_14, 
        p_wishbone_bd_ram_mem1_171_15, p_wishbone_bd_ram_mem1_172_8, 
        p_wishbone_bd_ram_mem1_172_9, p_wishbone_bd_ram_mem1_172_10, 
        p_wishbone_bd_ram_mem1_172_11, p_wishbone_bd_ram_mem1_172_12, 
        p_wishbone_bd_ram_mem1_172_13, p_wishbone_bd_ram_mem1_172_14, 
        p_wishbone_bd_ram_mem1_172_15, p_wishbone_bd_ram_mem1_173_8, 
        p_wishbone_bd_ram_mem1_173_9, p_wishbone_bd_ram_mem1_173_10, 
        p_wishbone_bd_ram_mem1_173_11, p_wishbone_bd_ram_mem1_173_12, 
        p_wishbone_bd_ram_mem1_173_13, p_wishbone_bd_ram_mem1_173_14, 
        p_wishbone_bd_ram_mem1_173_15, p_wishbone_bd_ram_mem1_174_8, 
        p_wishbone_bd_ram_mem1_174_9, p_wishbone_bd_ram_mem1_174_10, 
        p_wishbone_bd_ram_mem1_174_11, p_wishbone_bd_ram_mem1_174_12, 
        p_wishbone_bd_ram_mem1_174_13, p_wishbone_bd_ram_mem1_174_14, 
        p_wishbone_bd_ram_mem1_174_15, p_wishbone_bd_ram_mem1_175_8, 
        p_wishbone_bd_ram_mem1_175_9, p_wishbone_bd_ram_mem1_175_10, 
        p_wishbone_bd_ram_mem1_175_11, p_wishbone_bd_ram_mem1_175_12, 
        p_wishbone_bd_ram_mem1_175_13, p_wishbone_bd_ram_mem1_175_14, 
        p_wishbone_bd_ram_mem1_175_15, p_wishbone_bd_ram_mem1_176_8, 
        p_wishbone_bd_ram_mem1_176_9, p_wishbone_bd_ram_mem1_176_10, 
        p_wishbone_bd_ram_mem1_176_11, p_wishbone_bd_ram_mem1_176_12, 
        p_wishbone_bd_ram_mem1_176_13, p_wishbone_bd_ram_mem1_176_14, 
        p_wishbone_bd_ram_mem1_176_15, p_wishbone_bd_ram_mem1_177_8, 
        p_wishbone_bd_ram_mem1_177_9, p_wishbone_bd_ram_mem1_177_10, 
        p_wishbone_bd_ram_mem1_177_11, p_wishbone_bd_ram_mem1_177_12, 
        p_wishbone_bd_ram_mem1_177_13, p_wishbone_bd_ram_mem1_177_14, 
        p_wishbone_bd_ram_mem1_177_15, p_wishbone_bd_ram_mem1_178_8, 
        p_wishbone_bd_ram_mem1_178_9, p_wishbone_bd_ram_mem1_178_10, 
        p_wishbone_bd_ram_mem1_178_11, p_wishbone_bd_ram_mem1_178_12, 
        p_wishbone_bd_ram_mem1_178_13, p_wishbone_bd_ram_mem1_178_14, 
        p_wishbone_bd_ram_mem1_178_15, p_wishbone_bd_ram_mem1_179_8, 
        p_wishbone_bd_ram_mem1_179_9, p_wishbone_bd_ram_mem1_179_10, 
        p_wishbone_bd_ram_mem1_179_11, p_wishbone_bd_ram_mem1_179_12, 
        p_wishbone_bd_ram_mem1_179_13, p_wishbone_bd_ram_mem1_179_14, 
        p_wishbone_bd_ram_mem1_179_15, p_wishbone_bd_ram_mem1_180_8, 
        p_wishbone_bd_ram_mem1_180_9, p_wishbone_bd_ram_mem1_180_10, 
        p_wishbone_bd_ram_mem1_180_11, p_wishbone_bd_ram_mem1_180_12, 
        p_wishbone_bd_ram_mem1_180_13, p_wishbone_bd_ram_mem1_180_14, 
        p_wishbone_bd_ram_mem1_180_15, p_wishbone_bd_ram_mem1_181_8, 
        p_wishbone_bd_ram_mem1_181_9, p_wishbone_bd_ram_mem1_181_10, 
        p_wishbone_bd_ram_mem1_181_11, p_wishbone_bd_ram_mem1_181_12, 
        p_wishbone_bd_ram_mem1_181_13, p_wishbone_bd_ram_mem1_181_14, 
        p_wishbone_bd_ram_mem1_181_15, p_wishbone_bd_ram_mem1_182_8, 
        p_wishbone_bd_ram_mem1_182_9, p_wishbone_bd_ram_mem1_182_10, 
        p_wishbone_bd_ram_mem1_182_11, p_wishbone_bd_ram_mem1_182_12, 
        p_wishbone_bd_ram_mem1_182_13, p_wishbone_bd_ram_mem1_182_14, 
        p_wishbone_bd_ram_mem1_182_15, p_wishbone_bd_ram_mem1_183_8, 
        p_wishbone_bd_ram_mem1_183_9, p_wishbone_bd_ram_mem1_183_10, 
        p_wishbone_bd_ram_mem1_183_11, p_wishbone_bd_ram_mem1_183_12, 
        p_wishbone_bd_ram_mem1_183_13, p_wishbone_bd_ram_mem1_183_14, 
        p_wishbone_bd_ram_mem1_183_15, p_wishbone_bd_ram_mem1_184_8, 
        p_wishbone_bd_ram_mem1_184_9, p_wishbone_bd_ram_mem1_184_10, 
        p_wishbone_bd_ram_mem1_184_11, p_wishbone_bd_ram_mem1_184_12, 
        p_wishbone_bd_ram_mem1_184_13, p_wishbone_bd_ram_mem1_184_14, 
        p_wishbone_bd_ram_mem1_184_15, p_wishbone_bd_ram_mem1_185_8, 
        p_wishbone_bd_ram_mem1_185_9, p_wishbone_bd_ram_mem1_185_10, 
        p_wishbone_bd_ram_mem1_185_11, p_wishbone_bd_ram_mem1_185_12, 
        p_wishbone_bd_ram_mem1_185_13, p_wishbone_bd_ram_mem1_185_14, 
        p_wishbone_bd_ram_mem1_185_15, p_wishbone_bd_ram_mem1_186_8, 
        p_wishbone_bd_ram_mem1_186_9, p_wishbone_bd_ram_mem1_186_10, 
        p_wishbone_bd_ram_mem1_186_11, p_wishbone_bd_ram_mem1_186_12, 
        p_wishbone_bd_ram_mem1_186_13, p_wishbone_bd_ram_mem1_186_14, 
        p_wishbone_bd_ram_mem1_186_15, p_wishbone_bd_ram_mem1_187_8, 
        p_wishbone_bd_ram_mem1_187_9, p_wishbone_bd_ram_mem1_187_10, 
        p_wishbone_bd_ram_mem1_187_11, p_wishbone_bd_ram_mem1_187_12, 
        p_wishbone_bd_ram_mem1_187_13, p_wishbone_bd_ram_mem1_187_14, 
        p_wishbone_bd_ram_mem1_187_15, p_wishbone_bd_ram_mem1_188_8, 
        p_wishbone_bd_ram_mem1_188_9, p_wishbone_bd_ram_mem1_188_10, 
        p_wishbone_bd_ram_mem1_188_11, p_wishbone_bd_ram_mem1_188_12, 
        p_wishbone_bd_ram_mem1_188_13, p_wishbone_bd_ram_mem1_188_14, 
        p_wishbone_bd_ram_mem1_188_15, p_wishbone_bd_ram_mem1_189_8, 
        p_wishbone_bd_ram_mem1_189_9, p_wishbone_bd_ram_mem1_189_10, 
        p_wishbone_bd_ram_mem1_189_11, p_wishbone_bd_ram_mem1_189_12, 
        p_wishbone_bd_ram_mem1_189_13, p_wishbone_bd_ram_mem1_189_14, 
        p_wishbone_bd_ram_mem1_189_15, p_wishbone_bd_ram_mem1_190_8, 
        p_wishbone_bd_ram_mem1_190_9, p_wishbone_bd_ram_mem1_190_10, 
        p_wishbone_bd_ram_mem1_190_11, p_wishbone_bd_ram_mem1_190_12, 
        p_wishbone_bd_ram_mem1_190_13, p_wishbone_bd_ram_mem1_190_14, 
        p_wishbone_bd_ram_mem1_190_15, p_wishbone_bd_ram_mem1_191_8, 
        p_wishbone_bd_ram_mem1_191_9, p_wishbone_bd_ram_mem1_191_10, 
        p_wishbone_bd_ram_mem1_191_11, p_wishbone_bd_ram_mem1_191_12, 
        p_wishbone_bd_ram_mem1_191_13, p_wishbone_bd_ram_mem1_191_14, 
        p_wishbone_bd_ram_mem1_191_15, p_wishbone_bd_ram_mem1_192_8, 
        p_wishbone_bd_ram_mem1_192_9, p_wishbone_bd_ram_mem1_192_10, 
        p_wishbone_bd_ram_mem1_192_11, p_wishbone_bd_ram_mem1_192_12, 
        p_wishbone_bd_ram_mem1_192_13, p_wishbone_bd_ram_mem1_192_14, 
        p_wishbone_bd_ram_mem1_192_15, p_wishbone_bd_ram_mem1_193_8, 
        p_wishbone_bd_ram_mem1_193_9, p_wishbone_bd_ram_mem1_193_10, 
        p_wishbone_bd_ram_mem1_193_11, p_wishbone_bd_ram_mem1_193_12, 
        p_wishbone_bd_ram_mem1_193_13, p_wishbone_bd_ram_mem1_193_14, 
        p_wishbone_bd_ram_mem1_193_15, p_wishbone_bd_ram_mem1_194_8, 
        p_wishbone_bd_ram_mem1_194_9, p_wishbone_bd_ram_mem1_194_10, 
        p_wishbone_bd_ram_mem1_194_11, p_wishbone_bd_ram_mem1_194_12, 
        p_wishbone_bd_ram_mem1_194_13, p_wishbone_bd_ram_mem1_194_14, 
        p_wishbone_bd_ram_mem1_194_15, p_wishbone_bd_ram_mem1_195_8, 
        p_wishbone_bd_ram_mem1_195_9, p_wishbone_bd_ram_mem1_195_10, 
        p_wishbone_bd_ram_mem1_195_11, p_wishbone_bd_ram_mem1_195_12, 
        p_wishbone_bd_ram_mem1_195_13, p_wishbone_bd_ram_mem1_195_14, 
        p_wishbone_bd_ram_mem1_195_15, p_wishbone_bd_ram_mem1_196_8, 
        p_wishbone_bd_ram_mem1_196_9, p_wishbone_bd_ram_mem1_196_10, 
        p_wishbone_bd_ram_mem1_196_11, p_wishbone_bd_ram_mem1_196_12, 
        p_wishbone_bd_ram_mem1_196_13, p_wishbone_bd_ram_mem1_196_14, 
        p_wishbone_bd_ram_mem1_196_15, p_wishbone_bd_ram_mem1_197_8, 
        p_wishbone_bd_ram_mem1_197_9, p_wishbone_bd_ram_mem1_197_10, 
        p_wishbone_bd_ram_mem1_197_11, p_wishbone_bd_ram_mem1_197_12, 
        p_wishbone_bd_ram_mem1_197_13, p_wishbone_bd_ram_mem1_197_14, 
        p_wishbone_bd_ram_mem1_197_15, p_wishbone_bd_ram_mem1_198_8, 
        p_wishbone_bd_ram_mem1_198_9, p_wishbone_bd_ram_mem1_198_10, 
        p_wishbone_bd_ram_mem1_198_11, p_wishbone_bd_ram_mem1_198_12, 
        p_wishbone_bd_ram_mem1_198_13, p_wishbone_bd_ram_mem1_198_14, 
        p_wishbone_bd_ram_mem1_198_15, p_wishbone_bd_ram_mem1_199_8, 
        p_wishbone_bd_ram_mem1_199_9, p_wishbone_bd_ram_mem1_199_10, 
        p_wishbone_bd_ram_mem1_199_11, p_wishbone_bd_ram_mem1_199_12, 
        p_wishbone_bd_ram_mem1_199_13, p_wishbone_bd_ram_mem1_199_14, 
        p_wishbone_bd_ram_mem1_199_15, p_wishbone_bd_ram_mem1_200_8, 
        p_wishbone_bd_ram_mem1_200_9, p_wishbone_bd_ram_mem1_200_10, 
        p_wishbone_bd_ram_mem1_200_11, p_wishbone_bd_ram_mem1_200_12, 
        p_wishbone_bd_ram_mem1_200_13, p_wishbone_bd_ram_mem1_200_14, 
        p_wishbone_bd_ram_mem1_200_15, p_wishbone_bd_ram_mem1_201_8, 
        p_wishbone_bd_ram_mem1_201_9, p_wishbone_bd_ram_mem1_201_10, 
        p_wishbone_bd_ram_mem1_201_11, p_wishbone_bd_ram_mem1_201_12, 
        p_wishbone_bd_ram_mem1_201_13, p_wishbone_bd_ram_mem1_201_14, 
        p_wishbone_bd_ram_mem1_201_15, p_wishbone_bd_ram_mem1_202_8, 
        p_wishbone_bd_ram_mem1_202_9, p_wishbone_bd_ram_mem1_202_10, 
        p_wishbone_bd_ram_mem1_202_11, p_wishbone_bd_ram_mem1_202_12, 
        p_wishbone_bd_ram_mem1_202_13, p_wishbone_bd_ram_mem1_202_14, 
        p_wishbone_bd_ram_mem1_202_15, p_wishbone_bd_ram_mem1_203_8, 
        p_wishbone_bd_ram_mem1_203_9, p_wishbone_bd_ram_mem1_203_10, 
        p_wishbone_bd_ram_mem1_203_11, p_wishbone_bd_ram_mem1_203_12, 
        p_wishbone_bd_ram_mem1_203_13, p_wishbone_bd_ram_mem1_203_14, 
        p_wishbone_bd_ram_mem1_203_15, p_wishbone_bd_ram_mem1_204_8, 
        p_wishbone_bd_ram_mem1_204_9, p_wishbone_bd_ram_mem1_204_10, 
        p_wishbone_bd_ram_mem1_204_11, p_wishbone_bd_ram_mem1_204_12, 
        p_wishbone_bd_ram_mem1_204_13, p_wishbone_bd_ram_mem1_204_14, 
        p_wishbone_bd_ram_mem1_204_15, p_wishbone_bd_ram_mem1_205_8, 
        p_wishbone_bd_ram_mem1_205_9, p_wishbone_bd_ram_mem1_205_10, 
        p_wishbone_bd_ram_mem1_205_11, p_wishbone_bd_ram_mem1_205_12, 
        p_wishbone_bd_ram_mem1_205_13, p_wishbone_bd_ram_mem1_205_14, 
        p_wishbone_bd_ram_mem1_205_15, p_wishbone_bd_ram_mem1_206_8, 
        p_wishbone_bd_ram_mem1_206_9, p_wishbone_bd_ram_mem1_206_10, 
        p_wishbone_bd_ram_mem1_206_11, p_wishbone_bd_ram_mem1_206_12, 
        p_wishbone_bd_ram_mem1_206_13, p_wishbone_bd_ram_mem1_206_14, 
        p_wishbone_bd_ram_mem1_206_15, p_wishbone_bd_ram_mem1_207_8, 
        p_wishbone_bd_ram_mem1_207_9, p_wishbone_bd_ram_mem1_207_10, 
        p_wishbone_bd_ram_mem1_207_11, p_wishbone_bd_ram_mem1_207_12, 
        p_wishbone_bd_ram_mem1_207_13, p_wishbone_bd_ram_mem1_207_14, 
        p_wishbone_bd_ram_mem1_207_15, p_wishbone_bd_ram_mem1_208_8, 
        p_wishbone_bd_ram_mem1_208_9, p_wishbone_bd_ram_mem1_208_10, 
        p_wishbone_bd_ram_mem1_208_11, p_wishbone_bd_ram_mem1_208_12, 
        p_wishbone_bd_ram_mem1_208_13, p_wishbone_bd_ram_mem1_208_14, 
        p_wishbone_bd_ram_mem1_208_15, p_wishbone_bd_ram_mem1_209_8, 
        p_wishbone_bd_ram_mem1_209_9, p_wishbone_bd_ram_mem1_209_10, 
        p_wishbone_bd_ram_mem1_209_11, p_wishbone_bd_ram_mem1_209_12, 
        p_wishbone_bd_ram_mem1_209_13, p_wishbone_bd_ram_mem1_209_14, 
        p_wishbone_bd_ram_mem1_209_15, p_wishbone_bd_ram_mem1_210_8, 
        p_wishbone_bd_ram_mem1_210_9, p_wishbone_bd_ram_mem1_210_10, 
        p_wishbone_bd_ram_mem1_210_11, p_wishbone_bd_ram_mem1_210_12, 
        p_wishbone_bd_ram_mem1_210_13, p_wishbone_bd_ram_mem1_210_14, 
        p_wishbone_bd_ram_mem1_210_15, p_wishbone_bd_ram_mem1_211_8, 
        p_wishbone_bd_ram_mem1_211_9, p_wishbone_bd_ram_mem1_211_10, 
        p_wishbone_bd_ram_mem1_211_11, p_wishbone_bd_ram_mem1_211_12, 
        p_wishbone_bd_ram_mem1_211_13, p_wishbone_bd_ram_mem1_211_14, 
        p_wishbone_bd_ram_mem1_211_15, p_wishbone_bd_ram_mem1_212_8, 
        p_wishbone_bd_ram_mem1_212_9, p_wishbone_bd_ram_mem1_212_10, 
        p_wishbone_bd_ram_mem1_212_11, p_wishbone_bd_ram_mem1_212_12, 
        p_wishbone_bd_ram_mem1_212_13, p_wishbone_bd_ram_mem1_212_14, 
        p_wishbone_bd_ram_mem1_212_15, p_wishbone_bd_ram_mem1_213_8, 
        p_wishbone_bd_ram_mem1_213_9, p_wishbone_bd_ram_mem1_213_10, 
        p_wishbone_bd_ram_mem1_213_11, p_wishbone_bd_ram_mem1_213_12, 
        p_wishbone_bd_ram_mem1_213_13, p_wishbone_bd_ram_mem1_213_14, 
        p_wishbone_bd_ram_mem1_213_15, p_wishbone_bd_ram_mem1_214_8, 
        p_wishbone_bd_ram_mem1_214_9, p_wishbone_bd_ram_mem1_214_10, 
        p_wishbone_bd_ram_mem1_214_11, p_wishbone_bd_ram_mem1_214_12, 
        p_wishbone_bd_ram_mem1_214_13, p_wishbone_bd_ram_mem1_214_14, 
        p_wishbone_bd_ram_mem1_214_15, p_wishbone_bd_ram_mem1_215_8, 
        p_wishbone_bd_ram_mem1_215_9, p_wishbone_bd_ram_mem1_215_10, 
        p_wishbone_bd_ram_mem1_215_11, p_wishbone_bd_ram_mem1_215_12, 
        p_wishbone_bd_ram_mem1_215_13, p_wishbone_bd_ram_mem1_215_14, 
        p_wishbone_bd_ram_mem1_215_15, p_wishbone_bd_ram_mem1_216_8, 
        p_wishbone_bd_ram_mem1_216_9, p_wishbone_bd_ram_mem1_216_10, 
        p_wishbone_bd_ram_mem1_216_11, p_wishbone_bd_ram_mem1_216_12, 
        p_wishbone_bd_ram_mem1_216_13, p_wishbone_bd_ram_mem1_216_14, 
        p_wishbone_bd_ram_mem1_216_15, p_wishbone_bd_ram_mem1_217_8, 
        p_wishbone_bd_ram_mem1_217_9, p_wishbone_bd_ram_mem1_217_10, 
        p_wishbone_bd_ram_mem1_217_11, p_wishbone_bd_ram_mem1_217_12, 
        p_wishbone_bd_ram_mem1_217_13, p_wishbone_bd_ram_mem1_217_14, 
        p_wishbone_bd_ram_mem1_217_15, p_wishbone_bd_ram_mem1_218_8, 
        p_wishbone_bd_ram_mem1_218_9, p_wishbone_bd_ram_mem1_218_10, 
        p_wishbone_bd_ram_mem1_218_11, p_wishbone_bd_ram_mem1_218_12, 
        p_wishbone_bd_ram_mem1_218_13, p_wishbone_bd_ram_mem1_218_14, 
        p_wishbone_bd_ram_mem1_218_15, p_wishbone_bd_ram_mem1_219_8, 
        p_wishbone_bd_ram_mem1_219_9, p_wishbone_bd_ram_mem1_219_10, 
        p_wishbone_bd_ram_mem1_219_11, p_wishbone_bd_ram_mem1_219_12, 
        p_wishbone_bd_ram_mem1_219_13, p_wishbone_bd_ram_mem1_219_14, 
        p_wishbone_bd_ram_mem1_219_15, p_wishbone_bd_ram_mem1_220_8, 
        p_wishbone_bd_ram_mem1_220_9, p_wishbone_bd_ram_mem1_220_10, 
        p_wishbone_bd_ram_mem1_220_11, p_wishbone_bd_ram_mem1_220_12, 
        p_wishbone_bd_ram_mem1_220_13, p_wishbone_bd_ram_mem1_220_14, 
        p_wishbone_bd_ram_mem1_220_15, p_wishbone_bd_ram_mem1_221_8, 
        p_wishbone_bd_ram_mem1_221_9, p_wishbone_bd_ram_mem1_221_10, 
        p_wishbone_bd_ram_mem1_221_11, p_wishbone_bd_ram_mem1_221_12, 
        p_wishbone_bd_ram_mem1_221_13, p_wishbone_bd_ram_mem1_221_14, 
        p_wishbone_bd_ram_mem1_221_15, p_wishbone_bd_ram_mem1_222_8, 
        p_wishbone_bd_ram_mem1_222_9, p_wishbone_bd_ram_mem1_222_10, 
        p_wishbone_bd_ram_mem1_222_11, p_wishbone_bd_ram_mem1_222_12, 
        p_wishbone_bd_ram_mem1_222_13, p_wishbone_bd_ram_mem1_222_14, 
        p_wishbone_bd_ram_mem1_222_15, p_wishbone_bd_ram_mem1_223_8, 
        p_wishbone_bd_ram_mem1_223_9, p_wishbone_bd_ram_mem1_223_10, 
        p_wishbone_bd_ram_mem1_223_11, p_wishbone_bd_ram_mem1_223_12, 
        p_wishbone_bd_ram_mem1_223_13, p_wishbone_bd_ram_mem1_223_14, 
        p_wishbone_bd_ram_mem1_223_15, p_wishbone_bd_ram_mem1_224_8, 
        p_wishbone_bd_ram_mem1_224_9, p_wishbone_bd_ram_mem1_224_10, 
        p_wishbone_bd_ram_mem1_224_11, p_wishbone_bd_ram_mem1_224_12, 
        p_wishbone_bd_ram_mem1_224_13, p_wishbone_bd_ram_mem1_224_14, 
        p_wishbone_bd_ram_mem1_224_15, p_wishbone_bd_ram_mem1_225_8, 
        p_wishbone_bd_ram_mem1_225_9, p_wishbone_bd_ram_mem1_225_10, 
        p_wishbone_bd_ram_mem1_225_11, p_wishbone_bd_ram_mem1_225_12, 
        p_wishbone_bd_ram_mem1_225_13, p_wishbone_bd_ram_mem1_225_14, 
        p_wishbone_bd_ram_mem1_225_15, p_wishbone_bd_ram_mem1_226_8, 
        p_wishbone_bd_ram_mem1_226_9, p_wishbone_bd_ram_mem1_226_10, 
        p_wishbone_bd_ram_mem1_226_11, p_wishbone_bd_ram_mem1_226_12, 
        p_wishbone_bd_ram_mem1_226_13, p_wishbone_bd_ram_mem1_226_14, 
        p_wishbone_bd_ram_mem1_226_15, p_wishbone_bd_ram_mem1_227_8, 
        p_wishbone_bd_ram_mem1_227_9, p_wishbone_bd_ram_mem1_227_10, 
        p_wishbone_bd_ram_mem1_227_11, p_wishbone_bd_ram_mem1_227_12, 
        p_wishbone_bd_ram_mem1_227_13, p_wishbone_bd_ram_mem1_227_14, 
        p_wishbone_bd_ram_mem1_227_15, p_wishbone_bd_ram_mem1_228_8, 
        p_wishbone_bd_ram_mem1_228_9, p_wishbone_bd_ram_mem1_228_10, 
        p_wishbone_bd_ram_mem1_228_11, p_wishbone_bd_ram_mem1_228_12, 
        p_wishbone_bd_ram_mem1_228_13, p_wishbone_bd_ram_mem1_228_14, 
        p_wishbone_bd_ram_mem1_228_15, p_wishbone_bd_ram_mem1_229_8, 
        p_wishbone_bd_ram_mem1_229_9, p_wishbone_bd_ram_mem1_229_10, 
        p_wishbone_bd_ram_mem1_229_11, p_wishbone_bd_ram_mem1_229_12, 
        p_wishbone_bd_ram_mem1_229_13, p_wishbone_bd_ram_mem1_229_14, 
        p_wishbone_bd_ram_mem1_229_15, p_wishbone_bd_ram_mem1_230_8, 
        p_wishbone_bd_ram_mem1_230_9, p_wishbone_bd_ram_mem1_230_10, 
        p_wishbone_bd_ram_mem1_230_11, p_wishbone_bd_ram_mem1_230_12, 
        p_wishbone_bd_ram_mem1_230_13, p_wishbone_bd_ram_mem1_230_14, 
        p_wishbone_bd_ram_mem1_230_15, p_wishbone_bd_ram_mem1_231_8, 
        p_wishbone_bd_ram_mem1_231_9, p_wishbone_bd_ram_mem1_231_10, 
        p_wishbone_bd_ram_mem1_231_11, p_wishbone_bd_ram_mem1_231_12, 
        p_wishbone_bd_ram_mem1_231_13, p_wishbone_bd_ram_mem1_231_14, 
        p_wishbone_bd_ram_mem1_231_15, p_wishbone_bd_ram_mem1_232_8, 
        p_wishbone_bd_ram_mem1_232_9, p_wishbone_bd_ram_mem1_232_10, 
        p_wishbone_bd_ram_mem1_232_11, p_wishbone_bd_ram_mem1_232_12, 
        p_wishbone_bd_ram_mem1_232_13, p_wishbone_bd_ram_mem1_232_14, 
        p_wishbone_bd_ram_mem1_232_15, p_wishbone_bd_ram_mem1_233_8, 
        p_wishbone_bd_ram_mem1_233_9, p_wishbone_bd_ram_mem1_233_10, 
        p_wishbone_bd_ram_mem1_233_11, p_wishbone_bd_ram_mem1_233_12, 
        p_wishbone_bd_ram_mem1_233_13, p_wishbone_bd_ram_mem1_233_14, 
        p_wishbone_bd_ram_mem1_233_15, p_wishbone_bd_ram_mem1_234_8, 
        p_wishbone_bd_ram_mem1_234_9, p_wishbone_bd_ram_mem1_234_10, 
        p_wishbone_bd_ram_mem1_234_11, p_wishbone_bd_ram_mem1_234_12, 
        p_wishbone_bd_ram_mem1_234_13, p_wishbone_bd_ram_mem1_234_14, 
        p_wishbone_bd_ram_mem1_234_15, p_wishbone_bd_ram_mem1_235_8, 
        p_wishbone_bd_ram_mem1_235_9, p_wishbone_bd_ram_mem1_235_10, 
        p_wishbone_bd_ram_mem1_235_11, p_wishbone_bd_ram_mem1_235_12, 
        p_wishbone_bd_ram_mem1_235_13, p_wishbone_bd_ram_mem1_235_14, 
        p_wishbone_bd_ram_mem1_235_15, p_wishbone_bd_ram_mem1_236_8, 
        p_wishbone_bd_ram_mem1_236_9, p_wishbone_bd_ram_mem1_236_10, 
        p_wishbone_bd_ram_mem1_236_11, p_wishbone_bd_ram_mem1_236_12, 
        p_wishbone_bd_ram_mem1_236_13, p_wishbone_bd_ram_mem1_236_14, 
        p_wishbone_bd_ram_mem1_236_15, p_wishbone_bd_ram_mem1_237_8, 
        p_wishbone_bd_ram_mem1_237_9, p_wishbone_bd_ram_mem1_237_10, 
        p_wishbone_bd_ram_mem1_237_11, p_wishbone_bd_ram_mem1_237_12, 
        p_wishbone_bd_ram_mem1_237_13, p_wishbone_bd_ram_mem1_237_14, 
        p_wishbone_bd_ram_mem1_237_15, p_wishbone_bd_ram_mem1_238_8, 
        p_wishbone_bd_ram_mem1_238_9, p_wishbone_bd_ram_mem1_238_10, 
        p_wishbone_bd_ram_mem1_238_11, p_wishbone_bd_ram_mem1_238_12, 
        p_wishbone_bd_ram_mem1_238_13, p_wishbone_bd_ram_mem1_238_14, 
        p_wishbone_bd_ram_mem1_238_15, p_wishbone_bd_ram_mem1_239_8, 
        p_wishbone_bd_ram_mem1_239_9, p_wishbone_bd_ram_mem1_239_10, 
        p_wishbone_bd_ram_mem1_239_11, p_wishbone_bd_ram_mem1_239_12, 
        p_wishbone_bd_ram_mem1_239_13, p_wishbone_bd_ram_mem1_239_14, 
        p_wishbone_bd_ram_mem1_239_15, p_wishbone_bd_ram_mem1_240_8, 
        p_wishbone_bd_ram_mem1_240_9, p_wishbone_bd_ram_mem1_240_10, 
        p_wishbone_bd_ram_mem1_240_11, p_wishbone_bd_ram_mem1_240_12, 
        p_wishbone_bd_ram_mem1_240_13, p_wishbone_bd_ram_mem1_240_14, 
        p_wishbone_bd_ram_mem1_240_15, p_wishbone_bd_ram_mem1_241_8, 
        p_wishbone_bd_ram_mem1_241_9, p_wishbone_bd_ram_mem1_241_10, 
        p_wishbone_bd_ram_mem1_241_11, p_wishbone_bd_ram_mem1_241_12, 
        p_wishbone_bd_ram_mem1_241_13, p_wishbone_bd_ram_mem1_241_14, 
        p_wishbone_bd_ram_mem1_241_15, p_wishbone_bd_ram_mem1_242_8, 
        p_wishbone_bd_ram_mem1_242_9, p_wishbone_bd_ram_mem1_242_10, 
        p_wishbone_bd_ram_mem1_242_11, p_wishbone_bd_ram_mem1_242_12, 
        p_wishbone_bd_ram_mem1_242_13, p_wishbone_bd_ram_mem1_242_14, 
        p_wishbone_bd_ram_mem1_242_15, p_wishbone_bd_ram_mem1_243_8, 
        p_wishbone_bd_ram_mem1_243_9, p_wishbone_bd_ram_mem1_243_10, 
        p_wishbone_bd_ram_mem1_243_11, p_wishbone_bd_ram_mem1_243_12, 
        p_wishbone_bd_ram_mem1_243_13, p_wishbone_bd_ram_mem1_243_14, 
        p_wishbone_bd_ram_mem1_243_15, p_wishbone_bd_ram_mem1_244_8, 
        p_wishbone_bd_ram_mem1_244_9, p_wishbone_bd_ram_mem1_244_10, 
        p_wishbone_bd_ram_mem1_244_11, p_wishbone_bd_ram_mem1_244_12, 
        p_wishbone_bd_ram_mem1_244_13, p_wishbone_bd_ram_mem1_244_14, 
        p_wishbone_bd_ram_mem1_244_15, p_wishbone_bd_ram_mem1_245_8, 
        p_wishbone_bd_ram_mem1_245_9, p_wishbone_bd_ram_mem1_245_10, 
        p_wishbone_bd_ram_mem1_245_11, p_wishbone_bd_ram_mem1_245_12, 
        p_wishbone_bd_ram_mem1_245_13, p_wishbone_bd_ram_mem1_245_14, 
        p_wishbone_bd_ram_mem1_245_15, p_wishbone_bd_ram_mem1_246_8, 
        p_wishbone_bd_ram_mem1_246_9, p_wishbone_bd_ram_mem1_246_10, 
        p_wishbone_bd_ram_mem1_246_11, p_wishbone_bd_ram_mem1_246_12, 
        p_wishbone_bd_ram_mem1_246_13, p_wishbone_bd_ram_mem1_246_14, 
        p_wishbone_bd_ram_mem1_246_15, p_wishbone_bd_ram_mem1_247_8, 
        p_wishbone_bd_ram_mem1_247_9, p_wishbone_bd_ram_mem1_247_10, 
        p_wishbone_bd_ram_mem1_247_11, p_wishbone_bd_ram_mem1_247_12, 
        p_wishbone_bd_ram_mem1_247_13, p_wishbone_bd_ram_mem1_247_14, 
        p_wishbone_bd_ram_mem1_247_15, p_wishbone_bd_ram_mem1_248_8, 
        p_wishbone_bd_ram_mem1_248_9, p_wishbone_bd_ram_mem1_248_10, 
        p_wishbone_bd_ram_mem1_248_11, p_wishbone_bd_ram_mem1_248_12, 
        p_wishbone_bd_ram_mem1_248_13, p_wishbone_bd_ram_mem1_248_14, 
        p_wishbone_bd_ram_mem1_248_15, p_wishbone_bd_ram_mem1_249_8, 
        p_wishbone_bd_ram_mem1_249_9, p_wishbone_bd_ram_mem1_249_10, 
        p_wishbone_bd_ram_mem1_249_11, p_wishbone_bd_ram_mem1_249_12, 
        p_wishbone_bd_ram_mem1_249_13, p_wishbone_bd_ram_mem1_249_14, 
        p_wishbone_bd_ram_mem1_249_15, p_wishbone_bd_ram_mem1_250_8, 
        p_wishbone_bd_ram_mem1_250_9, p_wishbone_bd_ram_mem1_250_10, 
        p_wishbone_bd_ram_mem1_250_11, p_wishbone_bd_ram_mem1_250_12, 
        p_wishbone_bd_ram_mem1_250_13, p_wishbone_bd_ram_mem1_250_14, 
        p_wishbone_bd_ram_mem1_250_15, p_wishbone_bd_ram_mem1_251_8, 
        p_wishbone_bd_ram_mem1_251_9, p_wishbone_bd_ram_mem1_251_10, 
        p_wishbone_bd_ram_mem1_251_11, p_wishbone_bd_ram_mem1_251_12, 
        p_wishbone_bd_ram_mem1_251_13, p_wishbone_bd_ram_mem1_251_14, 
        p_wishbone_bd_ram_mem1_251_15, p_wishbone_bd_ram_mem1_252_8, 
        p_wishbone_bd_ram_mem1_252_9, p_wishbone_bd_ram_mem1_252_10, 
        p_wishbone_bd_ram_mem1_252_11, p_wishbone_bd_ram_mem1_252_12, 
        p_wishbone_bd_ram_mem1_252_13, p_wishbone_bd_ram_mem1_252_14, 
        p_wishbone_bd_ram_mem1_252_15, p_wishbone_bd_ram_mem1_253_8, 
        p_wishbone_bd_ram_mem1_253_9, p_wishbone_bd_ram_mem1_253_10, 
        p_wishbone_bd_ram_mem1_253_11, p_wishbone_bd_ram_mem1_253_12, 
        p_wishbone_bd_ram_mem1_253_13, p_wishbone_bd_ram_mem1_253_14, 
        p_wishbone_bd_ram_mem1_253_15, p_wishbone_bd_ram_mem1_254_8, 
        p_wishbone_bd_ram_mem1_254_9, p_wishbone_bd_ram_mem1_254_10, 
        p_wishbone_bd_ram_mem1_254_11, p_wishbone_bd_ram_mem1_254_12, 
        p_wishbone_bd_ram_mem1_254_13, p_wishbone_bd_ram_mem1_254_14, 
        p_wishbone_bd_ram_mem1_254_15, p_wishbone_bd_ram_mem1_255_8, 
        p_wishbone_bd_ram_mem1_255_9, p_wishbone_bd_ram_mem1_255_10, 
        p_wishbone_bd_ram_mem1_255_11, p_wishbone_bd_ram_mem1_255_12, 
        p_wishbone_bd_ram_mem1_255_13, p_wishbone_bd_ram_mem1_255_14, 
        p_wishbone_bd_ram_mem1_255_15, p_wishbone_bd_ram_mem0_0_0, 
        p_wishbone_bd_ram_mem0_0_1, p_wishbone_bd_ram_mem0_0_2, 
        p_wishbone_bd_ram_mem0_0_3, p_wishbone_bd_ram_mem0_0_4, 
        p_wishbone_bd_ram_mem0_0_5, p_wishbone_bd_ram_mem0_0_6, 
        p_wishbone_bd_ram_mem0_0_7, p_wishbone_bd_ram_mem0_1_0, 
        p_wishbone_bd_ram_mem0_1_1, p_wishbone_bd_ram_mem0_1_2, 
        p_wishbone_bd_ram_mem0_1_3, p_wishbone_bd_ram_mem0_1_4, 
        p_wishbone_bd_ram_mem0_1_5, p_wishbone_bd_ram_mem0_1_6, 
        p_wishbone_bd_ram_mem0_1_7, p_wishbone_bd_ram_mem0_2_0, 
        p_wishbone_bd_ram_mem0_2_1, p_wishbone_bd_ram_mem0_2_2, 
        p_wishbone_bd_ram_mem0_2_3, p_wishbone_bd_ram_mem0_2_4, 
        p_wishbone_bd_ram_mem0_2_5, p_wishbone_bd_ram_mem0_2_6, 
        p_wishbone_bd_ram_mem0_2_7, p_wishbone_bd_ram_mem0_3_0, 
        p_wishbone_bd_ram_mem0_3_1, p_wishbone_bd_ram_mem0_3_2, 
        p_wishbone_bd_ram_mem0_3_3, p_wishbone_bd_ram_mem0_3_4, 
        p_wishbone_bd_ram_mem0_3_5, p_wishbone_bd_ram_mem0_3_6, 
        p_wishbone_bd_ram_mem0_3_7, p_wishbone_bd_ram_mem0_4_0, 
        p_wishbone_bd_ram_mem0_4_1, p_wishbone_bd_ram_mem0_4_2, 
        p_wishbone_bd_ram_mem0_4_3, p_wishbone_bd_ram_mem0_4_4, 
        p_wishbone_bd_ram_mem0_4_5, p_wishbone_bd_ram_mem0_4_6, 
        p_wishbone_bd_ram_mem0_4_7, p_wishbone_bd_ram_mem0_5_0, 
        p_wishbone_bd_ram_mem0_5_1, p_wishbone_bd_ram_mem0_5_2, 
        p_wishbone_bd_ram_mem0_5_3, p_wishbone_bd_ram_mem0_5_4, 
        p_wishbone_bd_ram_mem0_5_5, p_wishbone_bd_ram_mem0_5_6, 
        p_wishbone_bd_ram_mem0_5_7, p_wishbone_bd_ram_mem0_6_0, 
        p_wishbone_bd_ram_mem0_6_1, p_wishbone_bd_ram_mem0_6_2, 
        p_wishbone_bd_ram_mem0_6_3, p_wishbone_bd_ram_mem0_6_4, 
        p_wishbone_bd_ram_mem0_6_5, p_wishbone_bd_ram_mem0_6_6, 
        p_wishbone_bd_ram_mem0_6_7, p_wishbone_bd_ram_mem0_7_0, 
        p_wishbone_bd_ram_mem0_7_1, p_wishbone_bd_ram_mem0_7_2, 
        p_wishbone_bd_ram_mem0_7_3, p_wishbone_bd_ram_mem0_7_4, 
        p_wishbone_bd_ram_mem0_7_5, p_wishbone_bd_ram_mem0_7_6, 
        p_wishbone_bd_ram_mem0_7_7, p_wishbone_bd_ram_mem0_8_0, 
        p_wishbone_bd_ram_mem0_8_1, p_wishbone_bd_ram_mem0_8_2, 
        p_wishbone_bd_ram_mem0_8_3, p_wishbone_bd_ram_mem0_8_4, 
        p_wishbone_bd_ram_mem0_8_5, p_wishbone_bd_ram_mem0_8_6, 
        p_wishbone_bd_ram_mem0_8_7, p_wishbone_bd_ram_mem0_9_0, 
        p_wishbone_bd_ram_mem0_9_1, p_wishbone_bd_ram_mem0_9_2, 
        p_wishbone_bd_ram_mem0_9_3, p_wishbone_bd_ram_mem0_9_4, 
        p_wishbone_bd_ram_mem0_9_5, p_wishbone_bd_ram_mem0_9_6, 
        p_wishbone_bd_ram_mem0_9_7, p_wishbone_bd_ram_mem0_10_0, 
        p_wishbone_bd_ram_mem0_10_1, p_wishbone_bd_ram_mem0_10_2, 
        p_wishbone_bd_ram_mem0_10_3, p_wishbone_bd_ram_mem0_10_4, 
        p_wishbone_bd_ram_mem0_10_5, p_wishbone_bd_ram_mem0_10_6, 
        p_wishbone_bd_ram_mem0_10_7, p_wishbone_bd_ram_mem0_11_0, 
        p_wishbone_bd_ram_mem0_11_1, p_wishbone_bd_ram_mem0_11_2, 
        p_wishbone_bd_ram_mem0_11_3, p_wishbone_bd_ram_mem0_11_4, 
        p_wishbone_bd_ram_mem0_11_5, p_wishbone_bd_ram_mem0_11_6, 
        p_wishbone_bd_ram_mem0_11_7, p_wishbone_bd_ram_mem0_12_0, 
        p_wishbone_bd_ram_mem0_12_1, p_wishbone_bd_ram_mem0_12_2, 
        p_wishbone_bd_ram_mem0_12_3, p_wishbone_bd_ram_mem0_12_4, 
        p_wishbone_bd_ram_mem0_12_5, p_wishbone_bd_ram_mem0_12_6, 
        p_wishbone_bd_ram_mem0_12_7, p_wishbone_bd_ram_mem0_13_0, 
        p_wishbone_bd_ram_mem0_13_1, p_wishbone_bd_ram_mem0_13_2, 
        p_wishbone_bd_ram_mem0_13_3, p_wishbone_bd_ram_mem0_13_4, 
        p_wishbone_bd_ram_mem0_13_5, p_wishbone_bd_ram_mem0_13_6, 
        p_wishbone_bd_ram_mem0_13_7, p_wishbone_bd_ram_mem0_14_0, 
        p_wishbone_bd_ram_mem0_14_1, p_wishbone_bd_ram_mem0_14_2, 
        p_wishbone_bd_ram_mem0_14_3, p_wishbone_bd_ram_mem0_14_4, 
        p_wishbone_bd_ram_mem0_14_5, p_wishbone_bd_ram_mem0_14_6, 
        p_wishbone_bd_ram_mem0_14_7, p_wishbone_bd_ram_mem0_15_0, 
        p_wishbone_bd_ram_mem0_15_1, p_wishbone_bd_ram_mem0_15_2, 
        p_wishbone_bd_ram_mem0_15_3, p_wishbone_bd_ram_mem0_15_4, 
        p_wishbone_bd_ram_mem0_15_5, p_wishbone_bd_ram_mem0_15_6, 
        p_wishbone_bd_ram_mem0_15_7, p_wishbone_bd_ram_mem0_16_0, 
        p_wishbone_bd_ram_mem0_16_1, p_wishbone_bd_ram_mem0_16_2, 
        p_wishbone_bd_ram_mem0_16_3, p_wishbone_bd_ram_mem0_16_4, 
        p_wishbone_bd_ram_mem0_16_5, p_wishbone_bd_ram_mem0_16_6, 
        p_wishbone_bd_ram_mem0_16_7, p_wishbone_bd_ram_mem0_17_0, 
        p_wishbone_bd_ram_mem0_17_1, p_wishbone_bd_ram_mem0_17_2, 
        p_wishbone_bd_ram_mem0_17_3, p_wishbone_bd_ram_mem0_17_4, 
        p_wishbone_bd_ram_mem0_17_5, p_wishbone_bd_ram_mem0_17_6, 
        p_wishbone_bd_ram_mem0_17_7, p_wishbone_bd_ram_mem0_18_0, 
        p_wishbone_bd_ram_mem0_18_1, p_wishbone_bd_ram_mem0_18_2, 
        p_wishbone_bd_ram_mem0_18_3, p_wishbone_bd_ram_mem0_18_4, 
        p_wishbone_bd_ram_mem0_18_5, p_wishbone_bd_ram_mem0_18_6, 
        p_wishbone_bd_ram_mem0_18_7, p_wishbone_bd_ram_mem0_19_0, 
        p_wishbone_bd_ram_mem0_19_1, p_wishbone_bd_ram_mem0_19_2, 
        p_wishbone_bd_ram_mem0_19_3, p_wishbone_bd_ram_mem0_19_4, 
        p_wishbone_bd_ram_mem0_19_5, p_wishbone_bd_ram_mem0_19_6, 
        p_wishbone_bd_ram_mem0_19_7, p_wishbone_bd_ram_mem0_20_0, 
        p_wishbone_bd_ram_mem0_20_1, p_wishbone_bd_ram_mem0_20_2, 
        p_wishbone_bd_ram_mem0_20_3, p_wishbone_bd_ram_mem0_20_4, 
        p_wishbone_bd_ram_mem0_20_5, p_wishbone_bd_ram_mem0_20_6, 
        p_wishbone_bd_ram_mem0_20_7, p_wishbone_bd_ram_mem0_21_0, 
        p_wishbone_bd_ram_mem0_21_1, p_wishbone_bd_ram_mem0_21_2, 
        p_wishbone_bd_ram_mem0_21_3, p_wishbone_bd_ram_mem0_21_4, 
        p_wishbone_bd_ram_mem0_21_5, p_wishbone_bd_ram_mem0_21_6, 
        p_wishbone_bd_ram_mem0_21_7, p_wishbone_bd_ram_mem0_22_0, 
        p_wishbone_bd_ram_mem0_22_1, p_wishbone_bd_ram_mem0_22_2, 
        p_wishbone_bd_ram_mem0_22_3, p_wishbone_bd_ram_mem0_22_4, 
        p_wishbone_bd_ram_mem0_22_5, p_wishbone_bd_ram_mem0_22_6, 
        p_wishbone_bd_ram_mem0_22_7, p_wishbone_bd_ram_mem0_23_0, 
        p_wishbone_bd_ram_mem0_23_1, p_wishbone_bd_ram_mem0_23_2, 
        p_wishbone_bd_ram_mem0_23_3, p_wishbone_bd_ram_mem0_23_4, 
        p_wishbone_bd_ram_mem0_23_5, p_wishbone_bd_ram_mem0_23_6, 
        p_wishbone_bd_ram_mem0_23_7, p_wishbone_bd_ram_mem0_24_0, 
        p_wishbone_bd_ram_mem0_24_1, p_wishbone_bd_ram_mem0_24_2, 
        p_wishbone_bd_ram_mem0_24_3, p_wishbone_bd_ram_mem0_24_4, 
        p_wishbone_bd_ram_mem0_24_5, p_wishbone_bd_ram_mem0_24_6, 
        p_wishbone_bd_ram_mem0_24_7, p_wishbone_bd_ram_mem0_25_0, 
        p_wishbone_bd_ram_mem0_25_1, p_wishbone_bd_ram_mem0_25_2, 
        p_wishbone_bd_ram_mem0_25_3, p_wishbone_bd_ram_mem0_25_4, 
        p_wishbone_bd_ram_mem0_25_5, p_wishbone_bd_ram_mem0_25_6, 
        p_wishbone_bd_ram_mem0_25_7, p_wishbone_bd_ram_mem0_26_0, 
        p_wishbone_bd_ram_mem0_26_1, p_wishbone_bd_ram_mem0_26_2, 
        p_wishbone_bd_ram_mem0_26_3, p_wishbone_bd_ram_mem0_26_4, 
        p_wishbone_bd_ram_mem0_26_5, p_wishbone_bd_ram_mem0_26_6, 
        p_wishbone_bd_ram_mem0_26_7, p_wishbone_bd_ram_mem0_27_0, 
        p_wishbone_bd_ram_mem0_27_1, p_wishbone_bd_ram_mem0_27_2, 
        p_wishbone_bd_ram_mem0_27_3, p_wishbone_bd_ram_mem0_27_4, 
        p_wishbone_bd_ram_mem0_27_5, p_wishbone_bd_ram_mem0_27_6, 
        p_wishbone_bd_ram_mem0_27_7, p_wishbone_bd_ram_mem0_28_0, 
        p_wishbone_bd_ram_mem0_28_1, p_wishbone_bd_ram_mem0_28_2, 
        p_wishbone_bd_ram_mem0_28_3, p_wishbone_bd_ram_mem0_28_4, 
        p_wishbone_bd_ram_mem0_28_5, p_wishbone_bd_ram_mem0_28_6, 
        p_wishbone_bd_ram_mem0_28_7, p_wishbone_bd_ram_mem0_29_0, 
        p_wishbone_bd_ram_mem0_29_1, p_wishbone_bd_ram_mem0_29_2, 
        p_wishbone_bd_ram_mem0_29_3, p_wishbone_bd_ram_mem0_29_4, 
        p_wishbone_bd_ram_mem0_29_5, p_wishbone_bd_ram_mem0_29_6, 
        p_wishbone_bd_ram_mem0_29_7, p_wishbone_bd_ram_mem0_30_0, 
        p_wishbone_bd_ram_mem0_30_1, p_wishbone_bd_ram_mem0_30_2, 
        p_wishbone_bd_ram_mem0_30_3, p_wishbone_bd_ram_mem0_30_4, 
        p_wishbone_bd_ram_mem0_30_5, p_wishbone_bd_ram_mem0_30_6, 
        p_wishbone_bd_ram_mem0_30_7, p_wishbone_bd_ram_mem0_31_0, 
        p_wishbone_bd_ram_mem0_31_1, p_wishbone_bd_ram_mem0_31_2, 
        p_wishbone_bd_ram_mem0_31_3, p_wishbone_bd_ram_mem0_31_4, 
        p_wishbone_bd_ram_mem0_31_5, p_wishbone_bd_ram_mem0_31_6, 
        p_wishbone_bd_ram_mem0_31_7, p_wishbone_bd_ram_mem0_32_0, 
        p_wishbone_bd_ram_mem0_32_1, p_wishbone_bd_ram_mem0_32_2, 
        p_wishbone_bd_ram_mem0_32_3, p_wishbone_bd_ram_mem0_32_4, 
        p_wishbone_bd_ram_mem0_32_5, p_wishbone_bd_ram_mem0_32_6, 
        p_wishbone_bd_ram_mem0_32_7, p_wishbone_bd_ram_mem0_33_0, 
        p_wishbone_bd_ram_mem0_33_1, p_wishbone_bd_ram_mem0_33_2, 
        p_wishbone_bd_ram_mem0_33_3, p_wishbone_bd_ram_mem0_33_4, 
        p_wishbone_bd_ram_mem0_33_5, p_wishbone_bd_ram_mem0_33_6, 
        p_wishbone_bd_ram_mem0_33_7, p_wishbone_bd_ram_mem0_34_0, 
        p_wishbone_bd_ram_mem0_34_1, p_wishbone_bd_ram_mem0_34_2, 
        p_wishbone_bd_ram_mem0_34_3, p_wishbone_bd_ram_mem0_34_4, 
        p_wishbone_bd_ram_mem0_34_5, p_wishbone_bd_ram_mem0_34_6, 
        p_wishbone_bd_ram_mem0_34_7, p_wishbone_bd_ram_mem0_35_0, 
        p_wishbone_bd_ram_mem0_35_1, p_wishbone_bd_ram_mem0_35_2, 
        p_wishbone_bd_ram_mem0_35_3, p_wishbone_bd_ram_mem0_35_4, 
        p_wishbone_bd_ram_mem0_35_5, p_wishbone_bd_ram_mem0_35_6, 
        p_wishbone_bd_ram_mem0_35_7, p_wishbone_bd_ram_mem0_36_0, 
        p_wishbone_bd_ram_mem0_36_1, p_wishbone_bd_ram_mem0_36_2, 
        p_wishbone_bd_ram_mem0_36_3, p_wishbone_bd_ram_mem0_36_4, 
        p_wishbone_bd_ram_mem0_36_5, p_wishbone_bd_ram_mem0_36_6, 
        p_wishbone_bd_ram_mem0_36_7, p_wishbone_bd_ram_mem0_37_0, 
        p_wishbone_bd_ram_mem0_37_1, p_wishbone_bd_ram_mem0_37_2, 
        p_wishbone_bd_ram_mem0_37_3, p_wishbone_bd_ram_mem0_37_4, 
        p_wishbone_bd_ram_mem0_37_5, p_wishbone_bd_ram_mem0_37_6, 
        p_wishbone_bd_ram_mem0_37_7, p_wishbone_bd_ram_mem0_38_0, 
        p_wishbone_bd_ram_mem0_38_1, p_wishbone_bd_ram_mem0_38_2, 
        p_wishbone_bd_ram_mem0_38_3, p_wishbone_bd_ram_mem0_38_4, 
        p_wishbone_bd_ram_mem0_38_5, p_wishbone_bd_ram_mem0_38_6, 
        p_wishbone_bd_ram_mem0_38_7, p_wishbone_bd_ram_mem0_39_0, 
        p_wishbone_bd_ram_mem0_39_1, p_wishbone_bd_ram_mem0_39_2, 
        p_wishbone_bd_ram_mem0_39_3, p_wishbone_bd_ram_mem0_39_4, 
        p_wishbone_bd_ram_mem0_39_5, p_wishbone_bd_ram_mem0_39_6, 
        p_wishbone_bd_ram_mem0_39_7, p_wishbone_bd_ram_mem0_40_0, 
        p_wishbone_bd_ram_mem0_40_1, p_wishbone_bd_ram_mem0_40_2, 
        p_wishbone_bd_ram_mem0_40_3, p_wishbone_bd_ram_mem0_40_4, 
        p_wishbone_bd_ram_mem0_40_5, p_wishbone_bd_ram_mem0_40_6, 
        p_wishbone_bd_ram_mem0_40_7, p_wishbone_bd_ram_mem0_41_0, 
        p_wishbone_bd_ram_mem0_41_1, p_wishbone_bd_ram_mem0_41_2, 
        p_wishbone_bd_ram_mem0_41_3, p_wishbone_bd_ram_mem0_41_4, 
        p_wishbone_bd_ram_mem0_41_5, p_wishbone_bd_ram_mem0_41_6, 
        p_wishbone_bd_ram_mem0_41_7, p_wishbone_bd_ram_mem0_42_0, 
        p_wishbone_bd_ram_mem0_42_1, p_wishbone_bd_ram_mem0_42_2, 
        p_wishbone_bd_ram_mem0_42_3, p_wishbone_bd_ram_mem0_42_4, 
        p_wishbone_bd_ram_mem0_42_5, p_wishbone_bd_ram_mem0_42_6, 
        p_wishbone_bd_ram_mem0_42_7, p_wishbone_bd_ram_mem0_43_0, 
        p_wishbone_bd_ram_mem0_43_1, p_wishbone_bd_ram_mem0_43_2, 
        p_wishbone_bd_ram_mem0_43_3, p_wishbone_bd_ram_mem0_43_4, 
        p_wishbone_bd_ram_mem0_43_5, p_wishbone_bd_ram_mem0_43_6, 
        p_wishbone_bd_ram_mem0_43_7, p_wishbone_bd_ram_mem0_44_0, 
        p_wishbone_bd_ram_mem0_44_1, p_wishbone_bd_ram_mem0_44_2, 
        p_wishbone_bd_ram_mem0_44_3, p_wishbone_bd_ram_mem0_44_4, 
        p_wishbone_bd_ram_mem0_44_5, p_wishbone_bd_ram_mem0_44_6, 
        p_wishbone_bd_ram_mem0_44_7, p_wishbone_bd_ram_mem0_45_0, 
        p_wishbone_bd_ram_mem0_45_1, p_wishbone_bd_ram_mem0_45_2, 
        p_wishbone_bd_ram_mem0_45_3, p_wishbone_bd_ram_mem0_45_4, 
        p_wishbone_bd_ram_mem0_45_5, p_wishbone_bd_ram_mem0_45_6, 
        p_wishbone_bd_ram_mem0_45_7, p_wishbone_bd_ram_mem0_46_0, 
        p_wishbone_bd_ram_mem0_46_1, p_wishbone_bd_ram_mem0_46_2, 
        p_wishbone_bd_ram_mem0_46_3, p_wishbone_bd_ram_mem0_46_4, 
        p_wishbone_bd_ram_mem0_46_5, p_wishbone_bd_ram_mem0_46_6, 
        p_wishbone_bd_ram_mem0_46_7, p_wishbone_bd_ram_mem0_47_0, 
        p_wishbone_bd_ram_mem0_47_1, p_wishbone_bd_ram_mem0_47_2, 
        p_wishbone_bd_ram_mem0_47_3, p_wishbone_bd_ram_mem0_47_4, 
        p_wishbone_bd_ram_mem0_47_5, p_wishbone_bd_ram_mem0_47_6, 
        p_wishbone_bd_ram_mem0_47_7, p_wishbone_bd_ram_mem0_48_0, 
        p_wishbone_bd_ram_mem0_48_1, p_wishbone_bd_ram_mem0_48_2, 
        p_wishbone_bd_ram_mem0_48_3, p_wishbone_bd_ram_mem0_48_4, 
        p_wishbone_bd_ram_mem0_48_5, p_wishbone_bd_ram_mem0_48_6, 
        p_wishbone_bd_ram_mem0_48_7, p_wishbone_bd_ram_mem0_49_0, 
        p_wishbone_bd_ram_mem0_49_1, p_wishbone_bd_ram_mem0_49_2, 
        p_wishbone_bd_ram_mem0_49_3, p_wishbone_bd_ram_mem0_49_4, 
        p_wishbone_bd_ram_mem0_49_5, p_wishbone_bd_ram_mem0_49_6, 
        p_wishbone_bd_ram_mem0_49_7, p_wishbone_bd_ram_mem0_50_0, 
        p_wishbone_bd_ram_mem0_50_1, p_wishbone_bd_ram_mem0_50_2, 
        p_wishbone_bd_ram_mem0_50_3, p_wishbone_bd_ram_mem0_50_4, 
        p_wishbone_bd_ram_mem0_50_5, p_wishbone_bd_ram_mem0_50_6, 
        p_wishbone_bd_ram_mem0_50_7, p_wishbone_bd_ram_mem0_51_0, 
        p_wishbone_bd_ram_mem0_51_1, p_wishbone_bd_ram_mem0_51_2, 
        p_wishbone_bd_ram_mem0_51_3, p_wishbone_bd_ram_mem0_51_4, 
        p_wishbone_bd_ram_mem0_51_5, p_wishbone_bd_ram_mem0_51_6, 
        p_wishbone_bd_ram_mem0_51_7, p_wishbone_bd_ram_mem0_52_0, 
        p_wishbone_bd_ram_mem0_52_1, p_wishbone_bd_ram_mem0_52_2, 
        p_wishbone_bd_ram_mem0_52_3, p_wishbone_bd_ram_mem0_52_4, 
        p_wishbone_bd_ram_mem0_52_5, p_wishbone_bd_ram_mem0_52_6, 
        p_wishbone_bd_ram_mem0_52_7, p_wishbone_bd_ram_mem0_53_0, 
        p_wishbone_bd_ram_mem0_53_1, p_wishbone_bd_ram_mem0_53_2, 
        p_wishbone_bd_ram_mem0_53_3, p_wishbone_bd_ram_mem0_53_4, 
        p_wishbone_bd_ram_mem0_53_5, p_wishbone_bd_ram_mem0_53_6, 
        p_wishbone_bd_ram_mem0_53_7, p_wishbone_bd_ram_mem0_54_0, 
        p_wishbone_bd_ram_mem0_54_1, p_wishbone_bd_ram_mem0_54_2, 
        p_wishbone_bd_ram_mem0_54_3, p_wishbone_bd_ram_mem0_54_4, 
        p_wishbone_bd_ram_mem0_54_5, p_wishbone_bd_ram_mem0_54_6, 
        p_wishbone_bd_ram_mem0_54_7, p_wishbone_bd_ram_mem0_55_0, 
        p_wishbone_bd_ram_mem0_55_1, p_wishbone_bd_ram_mem0_55_2, 
        p_wishbone_bd_ram_mem0_55_3, p_wishbone_bd_ram_mem0_55_4, 
        p_wishbone_bd_ram_mem0_55_5, p_wishbone_bd_ram_mem0_55_6, 
        p_wishbone_bd_ram_mem0_55_7, p_wishbone_bd_ram_mem0_56_0, 
        p_wishbone_bd_ram_mem0_56_1, p_wishbone_bd_ram_mem0_56_2, 
        p_wishbone_bd_ram_mem0_56_3, p_wishbone_bd_ram_mem0_56_4, 
        p_wishbone_bd_ram_mem0_56_5, p_wishbone_bd_ram_mem0_56_6, 
        p_wishbone_bd_ram_mem0_56_7, p_wishbone_bd_ram_mem0_57_0, 
        p_wishbone_bd_ram_mem0_57_1, p_wishbone_bd_ram_mem0_57_2, 
        p_wishbone_bd_ram_mem0_57_3, p_wishbone_bd_ram_mem0_57_4, 
        p_wishbone_bd_ram_mem0_57_5, p_wishbone_bd_ram_mem0_57_6, 
        p_wishbone_bd_ram_mem0_57_7, p_wishbone_bd_ram_mem0_58_0, 
        p_wishbone_bd_ram_mem0_58_1, p_wishbone_bd_ram_mem0_58_2, 
        p_wishbone_bd_ram_mem0_58_3, p_wishbone_bd_ram_mem0_58_4, 
        p_wishbone_bd_ram_mem0_58_5, p_wishbone_bd_ram_mem0_58_6, 
        p_wishbone_bd_ram_mem0_58_7, p_wishbone_bd_ram_mem0_59_0, 
        p_wishbone_bd_ram_mem0_59_1, p_wishbone_bd_ram_mem0_59_2, 
        p_wishbone_bd_ram_mem0_59_3, p_wishbone_bd_ram_mem0_59_4, 
        p_wishbone_bd_ram_mem0_59_5, p_wishbone_bd_ram_mem0_59_6, 
        p_wishbone_bd_ram_mem0_59_7, p_wishbone_bd_ram_mem0_60_0, 
        p_wishbone_bd_ram_mem0_60_1, p_wishbone_bd_ram_mem0_60_2, 
        p_wishbone_bd_ram_mem0_60_3, p_wishbone_bd_ram_mem0_60_4, 
        p_wishbone_bd_ram_mem0_60_5, p_wishbone_bd_ram_mem0_60_6, 
        p_wishbone_bd_ram_mem0_60_7, p_wishbone_bd_ram_mem0_61_0, 
        p_wishbone_bd_ram_mem0_61_1, p_wishbone_bd_ram_mem0_61_2, 
        p_wishbone_bd_ram_mem0_61_3, p_wishbone_bd_ram_mem0_61_4, 
        p_wishbone_bd_ram_mem0_61_5, p_wishbone_bd_ram_mem0_61_6, 
        p_wishbone_bd_ram_mem0_61_7, p_wishbone_bd_ram_mem0_62_0, 
        p_wishbone_bd_ram_mem0_62_1, p_wishbone_bd_ram_mem0_62_2, 
        p_wishbone_bd_ram_mem0_62_3, p_wishbone_bd_ram_mem0_62_4, 
        p_wishbone_bd_ram_mem0_62_5, p_wishbone_bd_ram_mem0_62_6, 
        p_wishbone_bd_ram_mem0_62_7, p_wishbone_bd_ram_mem0_63_0, 
        p_wishbone_bd_ram_mem0_63_1, p_wishbone_bd_ram_mem0_63_2, 
        p_wishbone_bd_ram_mem0_63_3, p_wishbone_bd_ram_mem0_63_4, 
        p_wishbone_bd_ram_mem0_63_5, p_wishbone_bd_ram_mem0_63_6, 
        p_wishbone_bd_ram_mem0_63_7, p_wishbone_bd_ram_mem0_64_0, 
        p_wishbone_bd_ram_mem0_64_1, p_wishbone_bd_ram_mem0_64_2, 
        p_wishbone_bd_ram_mem0_64_3, p_wishbone_bd_ram_mem0_64_4, 
        p_wishbone_bd_ram_mem0_64_5, p_wishbone_bd_ram_mem0_64_6, 
        p_wishbone_bd_ram_mem0_64_7, p_wishbone_bd_ram_mem0_65_0, 
        p_wishbone_bd_ram_mem0_65_1, p_wishbone_bd_ram_mem0_65_2, 
        p_wishbone_bd_ram_mem0_65_3, p_wishbone_bd_ram_mem0_65_4, 
        p_wishbone_bd_ram_mem0_65_5, p_wishbone_bd_ram_mem0_65_6, 
        p_wishbone_bd_ram_mem0_65_7, p_wishbone_bd_ram_mem0_66_0, 
        p_wishbone_bd_ram_mem0_66_1, p_wishbone_bd_ram_mem0_66_2, 
        p_wishbone_bd_ram_mem0_66_3, p_wishbone_bd_ram_mem0_66_4, 
        p_wishbone_bd_ram_mem0_66_5, p_wishbone_bd_ram_mem0_66_6, 
        p_wishbone_bd_ram_mem0_66_7, p_wishbone_bd_ram_mem0_67_0, 
        p_wishbone_bd_ram_mem0_67_1, p_wishbone_bd_ram_mem0_67_2, 
        p_wishbone_bd_ram_mem0_67_3, p_wishbone_bd_ram_mem0_67_4, 
        p_wishbone_bd_ram_mem0_67_5, p_wishbone_bd_ram_mem0_67_6, 
        p_wishbone_bd_ram_mem0_67_7, p_wishbone_bd_ram_mem0_68_0, 
        p_wishbone_bd_ram_mem0_68_1, p_wishbone_bd_ram_mem0_68_2, 
        p_wishbone_bd_ram_mem0_68_3, p_wishbone_bd_ram_mem0_68_4, 
        p_wishbone_bd_ram_mem0_68_5, p_wishbone_bd_ram_mem0_68_6, 
        p_wishbone_bd_ram_mem0_68_7, p_wishbone_bd_ram_mem0_69_0, 
        p_wishbone_bd_ram_mem0_69_1, p_wishbone_bd_ram_mem0_69_2, 
        p_wishbone_bd_ram_mem0_69_3, p_wishbone_bd_ram_mem0_69_4, 
        p_wishbone_bd_ram_mem0_69_5, p_wishbone_bd_ram_mem0_69_6, 
        p_wishbone_bd_ram_mem0_69_7, p_wishbone_bd_ram_mem0_70_0, 
        p_wishbone_bd_ram_mem0_70_1, p_wishbone_bd_ram_mem0_70_2, 
        p_wishbone_bd_ram_mem0_70_3, p_wishbone_bd_ram_mem0_70_4, 
        p_wishbone_bd_ram_mem0_70_5, p_wishbone_bd_ram_mem0_70_6, 
        p_wishbone_bd_ram_mem0_70_7, p_wishbone_bd_ram_mem0_71_0, 
        p_wishbone_bd_ram_mem0_71_1, p_wishbone_bd_ram_mem0_71_2, 
        p_wishbone_bd_ram_mem0_71_3, p_wishbone_bd_ram_mem0_71_4, 
        p_wishbone_bd_ram_mem0_71_5, p_wishbone_bd_ram_mem0_71_6, 
        p_wishbone_bd_ram_mem0_71_7, p_wishbone_bd_ram_mem0_72_0, 
        p_wishbone_bd_ram_mem0_72_1, p_wishbone_bd_ram_mem0_72_2, 
        p_wishbone_bd_ram_mem0_72_3, p_wishbone_bd_ram_mem0_72_4, 
        p_wishbone_bd_ram_mem0_72_5, p_wishbone_bd_ram_mem0_72_6, 
        p_wishbone_bd_ram_mem0_72_7, p_wishbone_bd_ram_mem0_73_0, 
        p_wishbone_bd_ram_mem0_73_1, p_wishbone_bd_ram_mem0_73_2, 
        p_wishbone_bd_ram_mem0_73_3, p_wishbone_bd_ram_mem0_73_4, 
        p_wishbone_bd_ram_mem0_73_5, p_wishbone_bd_ram_mem0_73_6, 
        p_wishbone_bd_ram_mem0_73_7, p_wishbone_bd_ram_mem0_74_0, 
        p_wishbone_bd_ram_mem0_74_1, p_wishbone_bd_ram_mem0_74_2, 
        p_wishbone_bd_ram_mem0_74_3, p_wishbone_bd_ram_mem0_74_4, 
        p_wishbone_bd_ram_mem0_74_5, p_wishbone_bd_ram_mem0_74_6, 
        p_wishbone_bd_ram_mem0_74_7, p_wishbone_bd_ram_mem0_75_0, 
        p_wishbone_bd_ram_mem0_75_1, p_wishbone_bd_ram_mem0_75_2, 
        p_wishbone_bd_ram_mem0_75_3, p_wishbone_bd_ram_mem0_75_4, 
        p_wishbone_bd_ram_mem0_75_5, p_wishbone_bd_ram_mem0_75_6, 
        p_wishbone_bd_ram_mem0_75_7, p_wishbone_bd_ram_mem0_76_0, 
        p_wishbone_bd_ram_mem0_76_1, p_wishbone_bd_ram_mem0_76_2, 
        p_wishbone_bd_ram_mem0_76_3, p_wishbone_bd_ram_mem0_76_4, 
        p_wishbone_bd_ram_mem0_76_5, p_wishbone_bd_ram_mem0_76_6, 
        p_wishbone_bd_ram_mem0_76_7, p_wishbone_bd_ram_mem0_77_0, 
        p_wishbone_bd_ram_mem0_77_1, p_wishbone_bd_ram_mem0_77_2, 
        p_wishbone_bd_ram_mem0_77_3, p_wishbone_bd_ram_mem0_77_4, 
        p_wishbone_bd_ram_mem0_77_5, p_wishbone_bd_ram_mem0_77_6, 
        p_wishbone_bd_ram_mem0_77_7, p_wishbone_bd_ram_mem0_78_0, 
        p_wishbone_bd_ram_mem0_78_1, p_wishbone_bd_ram_mem0_78_2, 
        p_wishbone_bd_ram_mem0_78_3, p_wishbone_bd_ram_mem0_78_4, 
        p_wishbone_bd_ram_mem0_78_5, p_wishbone_bd_ram_mem0_78_6, 
        p_wishbone_bd_ram_mem0_78_7, p_wishbone_bd_ram_mem0_79_0, 
        p_wishbone_bd_ram_mem0_79_1, p_wishbone_bd_ram_mem0_79_2, 
        p_wishbone_bd_ram_mem0_79_3, p_wishbone_bd_ram_mem0_79_4, 
        p_wishbone_bd_ram_mem0_79_5, p_wishbone_bd_ram_mem0_79_6, 
        p_wishbone_bd_ram_mem0_79_7, p_wishbone_bd_ram_mem0_80_0, 
        p_wishbone_bd_ram_mem0_80_1, p_wishbone_bd_ram_mem0_80_2, 
        p_wishbone_bd_ram_mem0_80_3, p_wishbone_bd_ram_mem0_80_4, 
        p_wishbone_bd_ram_mem0_80_5, p_wishbone_bd_ram_mem0_80_6, 
        p_wishbone_bd_ram_mem0_80_7, p_wishbone_bd_ram_mem0_81_0, 
        p_wishbone_bd_ram_mem0_81_1, p_wishbone_bd_ram_mem0_81_2, 
        p_wishbone_bd_ram_mem0_81_3, p_wishbone_bd_ram_mem0_81_4, 
        p_wishbone_bd_ram_mem0_81_5, p_wishbone_bd_ram_mem0_81_6, 
        p_wishbone_bd_ram_mem0_81_7, p_wishbone_bd_ram_mem0_82_0, 
        p_wishbone_bd_ram_mem0_82_1, p_wishbone_bd_ram_mem0_82_2, 
        p_wishbone_bd_ram_mem0_82_3, p_wishbone_bd_ram_mem0_82_4, 
        p_wishbone_bd_ram_mem0_82_5, p_wishbone_bd_ram_mem0_82_6, 
        p_wishbone_bd_ram_mem0_82_7, p_wishbone_bd_ram_mem0_83_0, 
        p_wishbone_bd_ram_mem0_83_1, p_wishbone_bd_ram_mem0_83_2, 
        p_wishbone_bd_ram_mem0_83_3, p_wishbone_bd_ram_mem0_83_4, 
        p_wishbone_bd_ram_mem0_83_5, p_wishbone_bd_ram_mem0_83_6, 
        p_wishbone_bd_ram_mem0_83_7, p_wishbone_bd_ram_mem0_84_0, 
        p_wishbone_bd_ram_mem0_84_1, p_wishbone_bd_ram_mem0_84_2, 
        p_wishbone_bd_ram_mem0_84_3, p_wishbone_bd_ram_mem0_84_4, 
        p_wishbone_bd_ram_mem0_84_5, p_wishbone_bd_ram_mem0_84_6, 
        p_wishbone_bd_ram_mem0_84_7, p_wishbone_bd_ram_mem0_85_0, 
        p_wishbone_bd_ram_mem0_85_1, p_wishbone_bd_ram_mem0_85_2, 
        p_wishbone_bd_ram_mem0_85_3, p_wishbone_bd_ram_mem0_85_4, 
        p_wishbone_bd_ram_mem0_85_5, p_wishbone_bd_ram_mem0_85_6, 
        p_wishbone_bd_ram_mem0_85_7, p_wishbone_bd_ram_mem0_86_0, 
        p_wishbone_bd_ram_mem0_86_1, p_wishbone_bd_ram_mem0_86_2, 
        p_wishbone_bd_ram_mem0_86_3, p_wishbone_bd_ram_mem0_86_4, 
        p_wishbone_bd_ram_mem0_86_5, p_wishbone_bd_ram_mem0_86_6, 
        p_wishbone_bd_ram_mem0_86_7, p_wishbone_bd_ram_mem0_87_0, 
        p_wishbone_bd_ram_mem0_87_1, p_wishbone_bd_ram_mem0_87_2, 
        p_wishbone_bd_ram_mem0_87_3, p_wishbone_bd_ram_mem0_87_4, 
        p_wishbone_bd_ram_mem0_87_5, p_wishbone_bd_ram_mem0_87_6, 
        p_wishbone_bd_ram_mem0_87_7, p_wishbone_bd_ram_mem0_88_0, 
        p_wishbone_bd_ram_mem0_88_1, p_wishbone_bd_ram_mem0_88_2, 
        p_wishbone_bd_ram_mem0_88_3, p_wishbone_bd_ram_mem0_88_4, 
        p_wishbone_bd_ram_mem0_88_5, p_wishbone_bd_ram_mem0_88_6, 
        p_wishbone_bd_ram_mem0_88_7, p_wishbone_bd_ram_mem0_89_0, 
        p_wishbone_bd_ram_mem0_89_1, p_wishbone_bd_ram_mem0_89_2, 
        p_wishbone_bd_ram_mem0_89_3, p_wishbone_bd_ram_mem0_89_4, 
        p_wishbone_bd_ram_mem0_89_5, p_wishbone_bd_ram_mem0_89_6, 
        p_wishbone_bd_ram_mem0_89_7, p_wishbone_bd_ram_mem0_90_0, 
        p_wishbone_bd_ram_mem0_90_1, p_wishbone_bd_ram_mem0_90_2, 
        p_wishbone_bd_ram_mem0_90_3, p_wishbone_bd_ram_mem0_90_4, 
        p_wishbone_bd_ram_mem0_90_5, p_wishbone_bd_ram_mem0_90_6, 
        p_wishbone_bd_ram_mem0_90_7, p_wishbone_bd_ram_mem0_91_0, 
        p_wishbone_bd_ram_mem0_91_1, p_wishbone_bd_ram_mem0_91_2, 
        p_wishbone_bd_ram_mem0_91_3, p_wishbone_bd_ram_mem0_91_4, 
        p_wishbone_bd_ram_mem0_91_5, p_wishbone_bd_ram_mem0_91_6, 
        p_wishbone_bd_ram_mem0_91_7, p_wishbone_bd_ram_mem0_92_0, 
        p_wishbone_bd_ram_mem0_92_1, p_wishbone_bd_ram_mem0_92_2, 
        p_wishbone_bd_ram_mem0_92_3, p_wishbone_bd_ram_mem0_92_4, 
        p_wishbone_bd_ram_mem0_92_5, p_wishbone_bd_ram_mem0_92_6, 
        p_wishbone_bd_ram_mem0_92_7, p_wishbone_bd_ram_mem0_93_0, 
        p_wishbone_bd_ram_mem0_93_1, p_wishbone_bd_ram_mem0_93_2, 
        p_wishbone_bd_ram_mem0_93_3, p_wishbone_bd_ram_mem0_93_4, 
        p_wishbone_bd_ram_mem0_93_5, p_wishbone_bd_ram_mem0_93_6, 
        p_wishbone_bd_ram_mem0_93_7, p_wishbone_bd_ram_mem0_94_0, 
        p_wishbone_bd_ram_mem0_94_1, p_wishbone_bd_ram_mem0_94_2, 
        p_wishbone_bd_ram_mem0_94_3, p_wishbone_bd_ram_mem0_94_4, 
        p_wishbone_bd_ram_mem0_94_5, p_wishbone_bd_ram_mem0_94_6, 
        p_wishbone_bd_ram_mem0_94_7, p_wishbone_bd_ram_mem0_95_0, 
        p_wishbone_bd_ram_mem0_95_1, p_wishbone_bd_ram_mem0_95_2, 
        p_wishbone_bd_ram_mem0_95_3, p_wishbone_bd_ram_mem0_95_4, 
        p_wishbone_bd_ram_mem0_95_5, p_wishbone_bd_ram_mem0_95_6, 
        p_wishbone_bd_ram_mem0_95_7, p_wishbone_bd_ram_mem0_96_0, 
        p_wishbone_bd_ram_mem0_96_1, p_wishbone_bd_ram_mem0_96_2, 
        p_wishbone_bd_ram_mem0_96_3, p_wishbone_bd_ram_mem0_96_4, 
        p_wishbone_bd_ram_mem0_96_5, p_wishbone_bd_ram_mem0_96_6, 
        p_wishbone_bd_ram_mem0_96_7, p_wishbone_bd_ram_mem0_97_0, 
        p_wishbone_bd_ram_mem0_97_1, p_wishbone_bd_ram_mem0_97_2, 
        p_wishbone_bd_ram_mem0_97_3, p_wishbone_bd_ram_mem0_97_4, 
        p_wishbone_bd_ram_mem0_97_5, p_wishbone_bd_ram_mem0_97_6, 
        p_wishbone_bd_ram_mem0_97_7, p_wishbone_bd_ram_mem0_98_0, 
        p_wishbone_bd_ram_mem0_98_1, p_wishbone_bd_ram_mem0_98_2, 
        p_wishbone_bd_ram_mem0_98_3, p_wishbone_bd_ram_mem0_98_4, 
        p_wishbone_bd_ram_mem0_98_5, p_wishbone_bd_ram_mem0_98_6, 
        p_wishbone_bd_ram_mem0_98_7, p_wishbone_bd_ram_mem0_99_0, 
        p_wishbone_bd_ram_mem0_99_1, p_wishbone_bd_ram_mem0_99_2, 
        p_wishbone_bd_ram_mem0_99_3, p_wishbone_bd_ram_mem0_99_4, 
        p_wishbone_bd_ram_mem0_99_5, p_wishbone_bd_ram_mem0_99_6, 
        p_wishbone_bd_ram_mem0_99_7, p_wishbone_bd_ram_mem0_100_0, 
        p_wishbone_bd_ram_mem0_100_1, p_wishbone_bd_ram_mem0_100_2, 
        p_wishbone_bd_ram_mem0_100_3, p_wishbone_bd_ram_mem0_100_4, 
        p_wishbone_bd_ram_mem0_100_5, p_wishbone_bd_ram_mem0_100_6, 
        p_wishbone_bd_ram_mem0_100_7, p_wishbone_bd_ram_mem0_101_0, 
        p_wishbone_bd_ram_mem0_101_1, p_wishbone_bd_ram_mem0_101_2, 
        p_wishbone_bd_ram_mem0_101_3, p_wishbone_bd_ram_mem0_101_4, 
        p_wishbone_bd_ram_mem0_101_5, p_wishbone_bd_ram_mem0_101_6, 
        p_wishbone_bd_ram_mem0_101_7, p_wishbone_bd_ram_mem0_102_0, 
        p_wishbone_bd_ram_mem0_102_1, p_wishbone_bd_ram_mem0_102_2, 
        p_wishbone_bd_ram_mem0_102_3, p_wishbone_bd_ram_mem0_102_4, 
        p_wishbone_bd_ram_mem0_102_5, p_wishbone_bd_ram_mem0_102_6, 
        p_wishbone_bd_ram_mem0_102_7, p_wishbone_bd_ram_mem0_103_0, 
        p_wishbone_bd_ram_mem0_103_1, p_wishbone_bd_ram_mem0_103_2, 
        p_wishbone_bd_ram_mem0_103_3, p_wishbone_bd_ram_mem0_103_4, 
        p_wishbone_bd_ram_mem0_103_5, p_wishbone_bd_ram_mem0_103_6, 
        p_wishbone_bd_ram_mem0_103_7, p_wishbone_bd_ram_mem0_104_0, 
        p_wishbone_bd_ram_mem0_104_1, p_wishbone_bd_ram_mem0_104_2, 
        p_wishbone_bd_ram_mem0_104_3, p_wishbone_bd_ram_mem0_104_4, 
        p_wishbone_bd_ram_mem0_104_5, p_wishbone_bd_ram_mem0_104_6, 
        p_wishbone_bd_ram_mem0_104_7, p_wishbone_bd_ram_mem0_105_0, 
        p_wishbone_bd_ram_mem0_105_1, p_wishbone_bd_ram_mem0_105_2, 
        p_wishbone_bd_ram_mem0_105_3, p_wishbone_bd_ram_mem0_105_4, 
        p_wishbone_bd_ram_mem0_105_5, p_wishbone_bd_ram_mem0_105_6, 
        p_wishbone_bd_ram_mem0_105_7, p_wishbone_bd_ram_mem0_106_0, 
        p_wishbone_bd_ram_mem0_106_1, p_wishbone_bd_ram_mem0_106_2, 
        p_wishbone_bd_ram_mem0_106_3, p_wishbone_bd_ram_mem0_106_4, 
        p_wishbone_bd_ram_mem0_106_5, p_wishbone_bd_ram_mem0_106_6, 
        p_wishbone_bd_ram_mem0_106_7, p_wishbone_bd_ram_mem0_107_0, 
        p_wishbone_bd_ram_mem0_107_1, p_wishbone_bd_ram_mem0_107_2, 
        p_wishbone_bd_ram_mem0_107_3, p_wishbone_bd_ram_mem0_107_4, 
        p_wishbone_bd_ram_mem0_107_5, p_wishbone_bd_ram_mem0_107_6, 
        p_wishbone_bd_ram_mem0_107_7, p_wishbone_bd_ram_mem0_108_0, 
        p_wishbone_bd_ram_mem0_108_1, p_wishbone_bd_ram_mem0_108_2, 
        p_wishbone_bd_ram_mem0_108_3, p_wishbone_bd_ram_mem0_108_4, 
        p_wishbone_bd_ram_mem0_108_5, p_wishbone_bd_ram_mem0_108_6, 
        p_wishbone_bd_ram_mem0_108_7, p_wishbone_bd_ram_mem0_109_0, 
        p_wishbone_bd_ram_mem0_109_1, p_wishbone_bd_ram_mem0_109_2, 
        p_wishbone_bd_ram_mem0_109_3, p_wishbone_bd_ram_mem0_109_4, 
        p_wishbone_bd_ram_mem0_109_5, p_wishbone_bd_ram_mem0_109_6, 
        p_wishbone_bd_ram_mem0_109_7, p_wishbone_bd_ram_mem0_110_0, 
        p_wishbone_bd_ram_mem0_110_1, p_wishbone_bd_ram_mem0_110_2, 
        p_wishbone_bd_ram_mem0_110_3, p_wishbone_bd_ram_mem0_110_4, 
        p_wishbone_bd_ram_mem0_110_5, p_wishbone_bd_ram_mem0_110_6, 
        p_wishbone_bd_ram_mem0_110_7, p_wishbone_bd_ram_mem0_111_0, 
        p_wishbone_bd_ram_mem0_111_1, p_wishbone_bd_ram_mem0_111_2, 
        p_wishbone_bd_ram_mem0_111_3, p_wishbone_bd_ram_mem0_111_4, 
        p_wishbone_bd_ram_mem0_111_5, p_wishbone_bd_ram_mem0_111_6, 
        p_wishbone_bd_ram_mem0_111_7, p_wishbone_bd_ram_mem0_112_0, 
        p_wishbone_bd_ram_mem0_112_1, p_wishbone_bd_ram_mem0_112_2, 
        p_wishbone_bd_ram_mem0_112_3, p_wishbone_bd_ram_mem0_112_4, 
        p_wishbone_bd_ram_mem0_112_5, p_wishbone_bd_ram_mem0_112_6, 
        p_wishbone_bd_ram_mem0_112_7, p_wishbone_bd_ram_mem0_113_0, 
        p_wishbone_bd_ram_mem0_113_1, p_wishbone_bd_ram_mem0_113_2, 
        p_wishbone_bd_ram_mem0_113_3, p_wishbone_bd_ram_mem0_113_4, 
        p_wishbone_bd_ram_mem0_113_5, p_wishbone_bd_ram_mem0_113_6, 
        p_wishbone_bd_ram_mem0_113_7, p_wishbone_bd_ram_mem0_114_0, 
        p_wishbone_bd_ram_mem0_114_1, p_wishbone_bd_ram_mem0_114_2, 
        p_wishbone_bd_ram_mem0_114_3, p_wishbone_bd_ram_mem0_114_4, 
        p_wishbone_bd_ram_mem0_114_5, p_wishbone_bd_ram_mem0_114_6, 
        p_wishbone_bd_ram_mem0_114_7, p_wishbone_bd_ram_mem0_115_0, 
        p_wishbone_bd_ram_mem0_115_1, p_wishbone_bd_ram_mem0_115_2, 
        p_wishbone_bd_ram_mem0_115_3, p_wishbone_bd_ram_mem0_115_4, 
        p_wishbone_bd_ram_mem0_115_5, p_wishbone_bd_ram_mem0_115_6, 
        p_wishbone_bd_ram_mem0_115_7, p_wishbone_bd_ram_mem0_116_0, 
        p_wishbone_bd_ram_mem0_116_1, p_wishbone_bd_ram_mem0_116_2, 
        p_wishbone_bd_ram_mem0_116_3, p_wishbone_bd_ram_mem0_116_4, 
        p_wishbone_bd_ram_mem0_116_5, p_wishbone_bd_ram_mem0_116_6, 
        p_wishbone_bd_ram_mem0_116_7, p_wishbone_bd_ram_mem0_117_0, 
        p_wishbone_bd_ram_mem0_117_1, p_wishbone_bd_ram_mem0_117_2, 
        p_wishbone_bd_ram_mem0_117_3, p_wishbone_bd_ram_mem0_117_4, 
        p_wishbone_bd_ram_mem0_117_5, p_wishbone_bd_ram_mem0_117_6, 
        p_wishbone_bd_ram_mem0_117_7, p_wishbone_bd_ram_mem0_118_0, 
        p_wishbone_bd_ram_mem0_118_1, p_wishbone_bd_ram_mem0_118_2, 
        p_wishbone_bd_ram_mem0_118_3, p_wishbone_bd_ram_mem0_118_4, 
        p_wishbone_bd_ram_mem0_118_5, p_wishbone_bd_ram_mem0_118_6, 
        p_wishbone_bd_ram_mem0_118_7, p_wishbone_bd_ram_mem0_119_0, 
        p_wishbone_bd_ram_mem0_119_1, p_wishbone_bd_ram_mem0_119_2, 
        p_wishbone_bd_ram_mem0_119_3, p_wishbone_bd_ram_mem0_119_4, 
        p_wishbone_bd_ram_mem0_119_5, p_wishbone_bd_ram_mem0_119_6, 
        p_wishbone_bd_ram_mem0_119_7, p_wishbone_bd_ram_mem0_120_0, 
        p_wishbone_bd_ram_mem0_120_1, p_wishbone_bd_ram_mem0_120_2, 
        p_wishbone_bd_ram_mem0_120_3, p_wishbone_bd_ram_mem0_120_4, 
        p_wishbone_bd_ram_mem0_120_5, p_wishbone_bd_ram_mem0_120_6, 
        p_wishbone_bd_ram_mem0_120_7, p_wishbone_bd_ram_mem0_121_0, 
        p_wishbone_bd_ram_mem0_121_1, p_wishbone_bd_ram_mem0_121_2, 
        p_wishbone_bd_ram_mem0_121_3, p_wishbone_bd_ram_mem0_121_4, 
        p_wishbone_bd_ram_mem0_121_5, p_wishbone_bd_ram_mem0_121_6, 
        p_wishbone_bd_ram_mem0_121_7, p_wishbone_bd_ram_mem0_122_0, 
        p_wishbone_bd_ram_mem0_122_1, p_wishbone_bd_ram_mem0_122_2, 
        p_wishbone_bd_ram_mem0_122_3, p_wishbone_bd_ram_mem0_122_4, 
        p_wishbone_bd_ram_mem0_122_5, p_wishbone_bd_ram_mem0_122_6, 
        p_wishbone_bd_ram_mem0_122_7, p_wishbone_bd_ram_mem0_123_0, 
        p_wishbone_bd_ram_mem0_123_1, p_wishbone_bd_ram_mem0_123_2, 
        p_wishbone_bd_ram_mem0_123_3, p_wishbone_bd_ram_mem0_123_4, 
        p_wishbone_bd_ram_mem0_123_5, p_wishbone_bd_ram_mem0_123_6, 
        p_wishbone_bd_ram_mem0_123_7, p_wishbone_bd_ram_mem0_124_0, 
        p_wishbone_bd_ram_mem0_124_1, p_wishbone_bd_ram_mem0_124_2, 
        p_wishbone_bd_ram_mem0_124_3, p_wishbone_bd_ram_mem0_124_4, 
        p_wishbone_bd_ram_mem0_124_5, p_wishbone_bd_ram_mem0_124_6, 
        p_wishbone_bd_ram_mem0_124_7, p_wishbone_bd_ram_mem0_125_0, 
        p_wishbone_bd_ram_mem0_125_1, p_wishbone_bd_ram_mem0_125_2, 
        p_wishbone_bd_ram_mem0_125_3, p_wishbone_bd_ram_mem0_125_4, 
        p_wishbone_bd_ram_mem0_125_5, p_wishbone_bd_ram_mem0_125_6, 
        p_wishbone_bd_ram_mem0_125_7, p_wishbone_bd_ram_mem0_126_0, 
        p_wishbone_bd_ram_mem0_126_1, p_wishbone_bd_ram_mem0_126_2, 
        p_wishbone_bd_ram_mem0_126_3, p_wishbone_bd_ram_mem0_126_4, 
        p_wishbone_bd_ram_mem0_126_5, p_wishbone_bd_ram_mem0_126_6, 
        p_wishbone_bd_ram_mem0_126_7, p_wishbone_bd_ram_mem0_127_0, 
        p_wishbone_bd_ram_mem0_127_1, p_wishbone_bd_ram_mem0_127_2, 
        p_wishbone_bd_ram_mem0_127_3, p_wishbone_bd_ram_mem0_127_4, 
        p_wishbone_bd_ram_mem0_127_5, p_wishbone_bd_ram_mem0_127_6, 
        p_wishbone_bd_ram_mem0_127_7, p_wishbone_bd_ram_mem0_128_0, 
        p_wishbone_bd_ram_mem0_128_1, p_wishbone_bd_ram_mem0_128_2, 
        p_wishbone_bd_ram_mem0_128_3, p_wishbone_bd_ram_mem0_128_4, 
        p_wishbone_bd_ram_mem0_128_5, p_wishbone_bd_ram_mem0_128_6, 
        p_wishbone_bd_ram_mem0_128_7, p_wishbone_bd_ram_mem0_129_0, 
        p_wishbone_bd_ram_mem0_129_1, p_wishbone_bd_ram_mem0_129_2, 
        p_wishbone_bd_ram_mem0_129_3, p_wishbone_bd_ram_mem0_129_4, 
        p_wishbone_bd_ram_mem0_129_5, p_wishbone_bd_ram_mem0_129_6, 
        p_wishbone_bd_ram_mem0_129_7, p_wishbone_bd_ram_mem0_130_0, 
        p_wishbone_bd_ram_mem0_130_1, p_wishbone_bd_ram_mem0_130_2, 
        p_wishbone_bd_ram_mem0_130_3, p_wishbone_bd_ram_mem0_130_4, 
        p_wishbone_bd_ram_mem0_130_5, p_wishbone_bd_ram_mem0_130_6, 
        p_wishbone_bd_ram_mem0_130_7, p_wishbone_bd_ram_mem0_131_0, 
        p_wishbone_bd_ram_mem0_131_1, p_wishbone_bd_ram_mem0_131_2, 
        p_wishbone_bd_ram_mem0_131_3, p_wishbone_bd_ram_mem0_131_4, 
        p_wishbone_bd_ram_mem0_131_5, p_wishbone_bd_ram_mem0_131_6, 
        p_wishbone_bd_ram_mem0_131_7, p_wishbone_bd_ram_mem0_132_0, 
        p_wishbone_bd_ram_mem0_132_1, p_wishbone_bd_ram_mem0_132_2, 
        p_wishbone_bd_ram_mem0_132_3, p_wishbone_bd_ram_mem0_132_4, 
        p_wishbone_bd_ram_mem0_132_5, p_wishbone_bd_ram_mem0_132_6, 
        p_wishbone_bd_ram_mem0_132_7, p_wishbone_bd_ram_mem0_133_0, 
        p_wishbone_bd_ram_mem0_133_1, p_wishbone_bd_ram_mem0_133_2, 
        p_wishbone_bd_ram_mem0_133_3, p_wishbone_bd_ram_mem0_133_4, 
        p_wishbone_bd_ram_mem0_133_5, p_wishbone_bd_ram_mem0_133_6, 
        p_wishbone_bd_ram_mem0_133_7, p_wishbone_bd_ram_mem0_134_0, 
        p_wishbone_bd_ram_mem0_134_1, p_wishbone_bd_ram_mem0_134_2, 
        p_wishbone_bd_ram_mem0_134_3, p_wishbone_bd_ram_mem0_134_4, 
        p_wishbone_bd_ram_mem0_134_5, p_wishbone_bd_ram_mem0_134_6, 
        p_wishbone_bd_ram_mem0_134_7, p_wishbone_bd_ram_mem0_135_0, 
        p_wishbone_bd_ram_mem0_135_1, p_wishbone_bd_ram_mem0_135_2, 
        p_wishbone_bd_ram_mem0_135_3, p_wishbone_bd_ram_mem0_135_4, 
        p_wishbone_bd_ram_mem0_135_5, p_wishbone_bd_ram_mem0_135_6, 
        p_wishbone_bd_ram_mem0_135_7, p_wishbone_bd_ram_mem0_136_0, 
        p_wishbone_bd_ram_mem0_136_1, p_wishbone_bd_ram_mem0_136_2, 
        p_wishbone_bd_ram_mem0_136_3, p_wishbone_bd_ram_mem0_136_4, 
        p_wishbone_bd_ram_mem0_136_5, p_wishbone_bd_ram_mem0_136_6, 
        p_wishbone_bd_ram_mem0_136_7, p_wishbone_bd_ram_mem0_137_0, 
        p_wishbone_bd_ram_mem0_137_1, p_wishbone_bd_ram_mem0_137_2, 
        p_wishbone_bd_ram_mem0_137_3, p_wishbone_bd_ram_mem0_137_4, 
        p_wishbone_bd_ram_mem0_137_5, p_wishbone_bd_ram_mem0_137_6, 
        p_wishbone_bd_ram_mem0_137_7, p_wishbone_bd_ram_mem0_138_0, 
        p_wishbone_bd_ram_mem0_138_1, p_wishbone_bd_ram_mem0_138_2, 
        p_wishbone_bd_ram_mem0_138_3, p_wishbone_bd_ram_mem0_138_4, 
        p_wishbone_bd_ram_mem0_138_5, p_wishbone_bd_ram_mem0_138_6, 
        p_wishbone_bd_ram_mem0_138_7, p_wishbone_bd_ram_mem0_139_0, 
        p_wishbone_bd_ram_mem0_139_1, p_wishbone_bd_ram_mem0_139_2, 
        p_wishbone_bd_ram_mem0_139_3, p_wishbone_bd_ram_mem0_139_4, 
        p_wishbone_bd_ram_mem0_139_5, p_wishbone_bd_ram_mem0_139_6, 
        p_wishbone_bd_ram_mem0_139_7, p_wishbone_bd_ram_mem0_140_0, 
        p_wishbone_bd_ram_mem0_140_1, p_wishbone_bd_ram_mem0_140_2, 
        p_wishbone_bd_ram_mem0_140_3, p_wishbone_bd_ram_mem0_140_4, 
        p_wishbone_bd_ram_mem0_140_5, p_wishbone_bd_ram_mem0_140_6, 
        p_wishbone_bd_ram_mem0_140_7, p_wishbone_bd_ram_mem0_141_0, 
        p_wishbone_bd_ram_mem0_141_1, p_wishbone_bd_ram_mem0_141_2, 
        p_wishbone_bd_ram_mem0_141_3, p_wishbone_bd_ram_mem0_141_4, 
        p_wishbone_bd_ram_mem0_141_5, p_wishbone_bd_ram_mem0_141_6, 
        p_wishbone_bd_ram_mem0_141_7, p_wishbone_bd_ram_mem0_142_0, 
        p_wishbone_bd_ram_mem0_142_1, p_wishbone_bd_ram_mem0_142_2, 
        p_wishbone_bd_ram_mem0_142_3, p_wishbone_bd_ram_mem0_142_4, 
        p_wishbone_bd_ram_mem0_142_5, p_wishbone_bd_ram_mem0_142_6, 
        p_wishbone_bd_ram_mem0_142_7, p_wishbone_bd_ram_mem0_143_0, 
        p_wishbone_bd_ram_mem0_143_1, p_wishbone_bd_ram_mem0_143_2, 
        p_wishbone_bd_ram_mem0_143_3, p_wishbone_bd_ram_mem0_143_4, 
        p_wishbone_bd_ram_mem0_143_5, p_wishbone_bd_ram_mem0_143_6, 
        p_wishbone_bd_ram_mem0_143_7, p_wishbone_bd_ram_mem0_144_0, 
        p_wishbone_bd_ram_mem0_144_1, p_wishbone_bd_ram_mem0_144_2, 
        p_wishbone_bd_ram_mem0_144_3, p_wishbone_bd_ram_mem0_144_4, 
        p_wishbone_bd_ram_mem0_144_5, p_wishbone_bd_ram_mem0_144_6, 
        p_wishbone_bd_ram_mem0_144_7, p_wishbone_bd_ram_mem0_145_0, 
        p_wishbone_bd_ram_mem0_145_1, p_wishbone_bd_ram_mem0_145_2, 
        p_wishbone_bd_ram_mem0_145_3, p_wishbone_bd_ram_mem0_145_4, 
        p_wishbone_bd_ram_mem0_145_5, p_wishbone_bd_ram_mem0_145_6, 
        p_wishbone_bd_ram_mem0_145_7, p_wishbone_bd_ram_mem0_146_0, 
        p_wishbone_bd_ram_mem0_146_1, p_wishbone_bd_ram_mem0_146_2, 
        p_wishbone_bd_ram_mem0_146_3, p_wishbone_bd_ram_mem0_146_4, 
        p_wishbone_bd_ram_mem0_146_5, p_wishbone_bd_ram_mem0_146_6, 
        p_wishbone_bd_ram_mem0_146_7, p_wishbone_bd_ram_mem0_147_0, 
        p_wishbone_bd_ram_mem0_147_1, p_wishbone_bd_ram_mem0_147_2, 
        p_wishbone_bd_ram_mem0_147_3, p_wishbone_bd_ram_mem0_147_4, 
        p_wishbone_bd_ram_mem0_147_5, p_wishbone_bd_ram_mem0_147_6, 
        p_wishbone_bd_ram_mem0_147_7, p_wishbone_bd_ram_mem0_148_0, 
        p_wishbone_bd_ram_mem0_148_1, p_wishbone_bd_ram_mem0_148_2, 
        p_wishbone_bd_ram_mem0_148_3, p_wishbone_bd_ram_mem0_148_4, 
        p_wishbone_bd_ram_mem0_148_5, p_wishbone_bd_ram_mem0_148_6, 
        p_wishbone_bd_ram_mem0_148_7, p_wishbone_bd_ram_mem0_149_0, 
        p_wishbone_bd_ram_mem0_149_1, p_wishbone_bd_ram_mem0_149_2, 
        p_wishbone_bd_ram_mem0_149_3, p_wishbone_bd_ram_mem0_149_4, 
        p_wishbone_bd_ram_mem0_149_5, p_wishbone_bd_ram_mem0_149_6, 
        p_wishbone_bd_ram_mem0_149_7, p_wishbone_bd_ram_mem0_150_0, 
        p_wishbone_bd_ram_mem0_150_1, p_wishbone_bd_ram_mem0_150_2, 
        p_wishbone_bd_ram_mem0_150_3, p_wishbone_bd_ram_mem0_150_4, 
        p_wishbone_bd_ram_mem0_150_5, p_wishbone_bd_ram_mem0_150_6, 
        p_wishbone_bd_ram_mem0_150_7, p_wishbone_bd_ram_mem0_151_0, 
        p_wishbone_bd_ram_mem0_151_1, p_wishbone_bd_ram_mem0_151_2, 
        p_wishbone_bd_ram_mem0_151_3, p_wishbone_bd_ram_mem0_151_4, 
        p_wishbone_bd_ram_mem0_151_5, p_wishbone_bd_ram_mem0_151_6, 
        p_wishbone_bd_ram_mem0_151_7, p_wishbone_bd_ram_mem0_152_0, 
        p_wishbone_bd_ram_mem0_152_1, p_wishbone_bd_ram_mem0_152_2, 
        p_wishbone_bd_ram_mem0_152_3, p_wishbone_bd_ram_mem0_152_4, 
        p_wishbone_bd_ram_mem0_152_5, p_wishbone_bd_ram_mem0_152_6, 
        p_wishbone_bd_ram_mem0_152_7, p_wishbone_bd_ram_mem0_153_0, 
        p_wishbone_bd_ram_mem0_153_1, p_wishbone_bd_ram_mem0_153_2, 
        p_wishbone_bd_ram_mem0_153_3, p_wishbone_bd_ram_mem0_153_4, 
        p_wishbone_bd_ram_mem0_153_5, p_wishbone_bd_ram_mem0_153_6, 
        p_wishbone_bd_ram_mem0_153_7, p_wishbone_bd_ram_mem0_154_0, 
        p_wishbone_bd_ram_mem0_154_1, p_wishbone_bd_ram_mem0_154_2, 
        p_wishbone_bd_ram_mem0_154_3, p_wishbone_bd_ram_mem0_154_4, 
        p_wishbone_bd_ram_mem0_154_5, p_wishbone_bd_ram_mem0_154_6, 
        p_wishbone_bd_ram_mem0_154_7, p_wishbone_bd_ram_mem0_155_0, 
        p_wishbone_bd_ram_mem0_155_1, p_wishbone_bd_ram_mem0_155_2, 
        p_wishbone_bd_ram_mem0_155_3, p_wishbone_bd_ram_mem0_155_4, 
        p_wishbone_bd_ram_mem0_155_5, p_wishbone_bd_ram_mem0_155_6, 
        p_wishbone_bd_ram_mem0_155_7, p_wishbone_bd_ram_mem0_156_0, 
        p_wishbone_bd_ram_mem0_156_1, p_wishbone_bd_ram_mem0_156_2, 
        p_wishbone_bd_ram_mem0_156_3, p_wishbone_bd_ram_mem0_156_4, 
        p_wishbone_bd_ram_mem0_156_5, p_wishbone_bd_ram_mem0_156_6, 
        p_wishbone_bd_ram_mem0_156_7, p_wishbone_bd_ram_mem0_157_0, 
        p_wishbone_bd_ram_mem0_157_1, p_wishbone_bd_ram_mem0_157_2, 
        p_wishbone_bd_ram_mem0_157_3, p_wishbone_bd_ram_mem0_157_4, 
        p_wishbone_bd_ram_mem0_157_5, p_wishbone_bd_ram_mem0_157_6, 
        p_wishbone_bd_ram_mem0_157_7, p_wishbone_bd_ram_mem0_158_0, 
        p_wishbone_bd_ram_mem0_158_1, p_wishbone_bd_ram_mem0_158_2, 
        p_wishbone_bd_ram_mem0_158_3, p_wishbone_bd_ram_mem0_158_4, 
        p_wishbone_bd_ram_mem0_158_5, p_wishbone_bd_ram_mem0_158_6, 
        p_wishbone_bd_ram_mem0_158_7, p_wishbone_bd_ram_mem0_159_0, 
        p_wishbone_bd_ram_mem0_159_1, p_wishbone_bd_ram_mem0_159_2, 
        p_wishbone_bd_ram_mem0_159_3, p_wishbone_bd_ram_mem0_159_4, 
        p_wishbone_bd_ram_mem0_159_5, p_wishbone_bd_ram_mem0_159_6, 
        p_wishbone_bd_ram_mem0_159_7, p_wishbone_bd_ram_mem0_160_0, 
        p_wishbone_bd_ram_mem0_160_1, p_wishbone_bd_ram_mem0_160_2, 
        p_wishbone_bd_ram_mem0_160_3, p_wishbone_bd_ram_mem0_160_4, 
        p_wishbone_bd_ram_mem0_160_5, p_wishbone_bd_ram_mem0_160_6, 
        p_wishbone_bd_ram_mem0_160_7, p_wishbone_bd_ram_mem0_161_0, 
        p_wishbone_bd_ram_mem0_161_1, p_wishbone_bd_ram_mem0_161_2, 
        p_wishbone_bd_ram_mem0_161_3, p_wishbone_bd_ram_mem0_161_4, 
        p_wishbone_bd_ram_mem0_161_5, p_wishbone_bd_ram_mem0_161_6, 
        p_wishbone_bd_ram_mem0_161_7, p_wishbone_bd_ram_mem0_162_0, 
        p_wishbone_bd_ram_mem0_162_1, p_wishbone_bd_ram_mem0_162_2, 
        p_wishbone_bd_ram_mem0_162_3, p_wishbone_bd_ram_mem0_162_4, 
        p_wishbone_bd_ram_mem0_162_5, p_wishbone_bd_ram_mem0_162_6, 
        p_wishbone_bd_ram_mem0_162_7, p_wishbone_bd_ram_mem0_163_0, 
        p_wishbone_bd_ram_mem0_163_1, p_wishbone_bd_ram_mem0_163_2, 
        p_wishbone_bd_ram_mem0_163_3, p_wishbone_bd_ram_mem0_163_4, 
        p_wishbone_bd_ram_mem0_163_5, p_wishbone_bd_ram_mem0_163_6, 
        p_wishbone_bd_ram_mem0_163_7, p_wishbone_bd_ram_mem0_164_0, 
        p_wishbone_bd_ram_mem0_164_1, p_wishbone_bd_ram_mem0_164_2, 
        p_wishbone_bd_ram_mem0_164_3, p_wishbone_bd_ram_mem0_164_4, 
        p_wishbone_bd_ram_mem0_164_5, p_wishbone_bd_ram_mem0_164_6, 
        p_wishbone_bd_ram_mem0_164_7, p_wishbone_bd_ram_mem0_165_0, 
        p_wishbone_bd_ram_mem0_165_1, p_wishbone_bd_ram_mem0_165_2, 
        p_wishbone_bd_ram_mem0_165_3, p_wishbone_bd_ram_mem0_165_4, 
        p_wishbone_bd_ram_mem0_165_5, p_wishbone_bd_ram_mem0_165_6, 
        p_wishbone_bd_ram_mem0_165_7, p_wishbone_bd_ram_mem0_166_0, 
        p_wishbone_bd_ram_mem0_166_1, p_wishbone_bd_ram_mem0_166_2, 
        p_wishbone_bd_ram_mem0_166_3, p_wishbone_bd_ram_mem0_166_4, 
        p_wishbone_bd_ram_mem0_166_5, p_wishbone_bd_ram_mem0_166_6, 
        p_wishbone_bd_ram_mem0_166_7, p_wishbone_bd_ram_mem0_167_0, 
        p_wishbone_bd_ram_mem0_167_1, p_wishbone_bd_ram_mem0_167_2, 
        p_wishbone_bd_ram_mem0_167_3, p_wishbone_bd_ram_mem0_167_4, 
        p_wishbone_bd_ram_mem0_167_5, p_wishbone_bd_ram_mem0_167_6, 
        p_wishbone_bd_ram_mem0_167_7, p_wishbone_bd_ram_mem0_168_0, 
        p_wishbone_bd_ram_mem0_168_1, p_wishbone_bd_ram_mem0_168_2, 
        p_wishbone_bd_ram_mem0_168_3, p_wishbone_bd_ram_mem0_168_4, 
        p_wishbone_bd_ram_mem0_168_5, p_wishbone_bd_ram_mem0_168_6, 
        p_wishbone_bd_ram_mem0_168_7, p_wishbone_bd_ram_mem0_169_0, 
        p_wishbone_bd_ram_mem0_169_1, p_wishbone_bd_ram_mem0_169_2, 
        p_wishbone_bd_ram_mem0_169_3, p_wishbone_bd_ram_mem0_169_4, 
        p_wishbone_bd_ram_mem0_169_5, p_wishbone_bd_ram_mem0_169_6, 
        p_wishbone_bd_ram_mem0_169_7, p_wishbone_bd_ram_mem0_170_0, 
        p_wishbone_bd_ram_mem0_170_1, p_wishbone_bd_ram_mem0_170_2, 
        p_wishbone_bd_ram_mem0_170_3, p_wishbone_bd_ram_mem0_170_4, 
        p_wishbone_bd_ram_mem0_170_5, p_wishbone_bd_ram_mem0_170_6, 
        p_wishbone_bd_ram_mem0_170_7, p_wishbone_bd_ram_mem0_171_0, 
        p_wishbone_bd_ram_mem0_171_1, p_wishbone_bd_ram_mem0_171_2, 
        p_wishbone_bd_ram_mem0_171_3, p_wishbone_bd_ram_mem0_171_4, 
        p_wishbone_bd_ram_mem0_171_5, p_wishbone_bd_ram_mem0_171_6, 
        p_wishbone_bd_ram_mem0_171_7, p_wishbone_bd_ram_mem0_172_0, 
        p_wishbone_bd_ram_mem0_172_1, p_wishbone_bd_ram_mem0_172_2, 
        p_wishbone_bd_ram_mem0_172_3, p_wishbone_bd_ram_mem0_172_4, 
        p_wishbone_bd_ram_mem0_172_5, p_wishbone_bd_ram_mem0_172_6, 
        p_wishbone_bd_ram_mem0_172_7, p_wishbone_bd_ram_mem0_173_0, 
        p_wishbone_bd_ram_mem0_173_1, p_wishbone_bd_ram_mem0_173_2, 
        p_wishbone_bd_ram_mem0_173_3, p_wishbone_bd_ram_mem0_173_4, 
        p_wishbone_bd_ram_mem0_173_5, p_wishbone_bd_ram_mem0_173_6, 
        p_wishbone_bd_ram_mem0_173_7, p_wishbone_bd_ram_mem0_174_0, 
        p_wishbone_bd_ram_mem0_174_1, p_wishbone_bd_ram_mem0_174_2, 
        p_wishbone_bd_ram_mem0_174_3, p_wishbone_bd_ram_mem0_174_4, 
        p_wishbone_bd_ram_mem0_174_5, p_wishbone_bd_ram_mem0_174_6, 
        p_wishbone_bd_ram_mem0_174_7, p_wishbone_bd_ram_mem0_175_0, 
        p_wishbone_bd_ram_mem0_175_1, p_wishbone_bd_ram_mem0_175_2, 
        p_wishbone_bd_ram_mem0_175_3, p_wishbone_bd_ram_mem0_175_4, 
        p_wishbone_bd_ram_mem0_175_5, p_wishbone_bd_ram_mem0_175_6, 
        p_wishbone_bd_ram_mem0_175_7, p_wishbone_bd_ram_mem0_176_0, 
        p_wishbone_bd_ram_mem0_176_1, p_wishbone_bd_ram_mem0_176_2, 
        p_wishbone_bd_ram_mem0_176_3, p_wishbone_bd_ram_mem0_176_4, 
        p_wishbone_bd_ram_mem0_176_5, p_wishbone_bd_ram_mem0_176_6, 
        p_wishbone_bd_ram_mem0_176_7, p_wishbone_bd_ram_mem0_177_0, 
        p_wishbone_bd_ram_mem0_177_1, p_wishbone_bd_ram_mem0_177_2, 
        p_wishbone_bd_ram_mem0_177_3, p_wishbone_bd_ram_mem0_177_4, 
        p_wishbone_bd_ram_mem0_177_5, p_wishbone_bd_ram_mem0_177_6, 
        p_wishbone_bd_ram_mem0_177_7, p_wishbone_bd_ram_mem0_178_0, 
        p_wishbone_bd_ram_mem0_178_1, p_wishbone_bd_ram_mem0_178_2, 
        p_wishbone_bd_ram_mem0_178_3, p_wishbone_bd_ram_mem0_178_4, 
        p_wishbone_bd_ram_mem0_178_5, p_wishbone_bd_ram_mem0_178_6, 
        p_wishbone_bd_ram_mem0_178_7, p_wishbone_bd_ram_mem0_179_0, 
        p_wishbone_bd_ram_mem0_179_1, p_wishbone_bd_ram_mem0_179_2, 
        p_wishbone_bd_ram_mem0_179_3, p_wishbone_bd_ram_mem0_179_4, 
        p_wishbone_bd_ram_mem0_179_5, p_wishbone_bd_ram_mem0_179_6, 
        p_wishbone_bd_ram_mem0_179_7, p_wishbone_bd_ram_mem0_180_0, 
        p_wishbone_bd_ram_mem0_180_1, p_wishbone_bd_ram_mem0_180_2, 
        p_wishbone_bd_ram_mem0_180_3, p_wishbone_bd_ram_mem0_180_4, 
        p_wishbone_bd_ram_mem0_180_5, p_wishbone_bd_ram_mem0_180_6, 
        p_wishbone_bd_ram_mem0_180_7, p_wishbone_bd_ram_mem0_181_0, 
        p_wishbone_bd_ram_mem0_181_1, p_wishbone_bd_ram_mem0_181_2, 
        p_wishbone_bd_ram_mem0_181_3, p_wishbone_bd_ram_mem0_181_4, 
        p_wishbone_bd_ram_mem0_181_5, p_wishbone_bd_ram_mem0_181_6, 
        p_wishbone_bd_ram_mem0_181_7, p_wishbone_bd_ram_mem0_182_0, 
        p_wishbone_bd_ram_mem0_182_1, p_wishbone_bd_ram_mem0_182_2, 
        p_wishbone_bd_ram_mem0_182_3, p_wishbone_bd_ram_mem0_182_4, 
        p_wishbone_bd_ram_mem0_182_5, p_wishbone_bd_ram_mem0_182_6, 
        p_wishbone_bd_ram_mem0_182_7, p_wishbone_bd_ram_mem0_183_0, 
        p_wishbone_bd_ram_mem0_183_1, p_wishbone_bd_ram_mem0_183_2, 
        p_wishbone_bd_ram_mem0_183_3, p_wishbone_bd_ram_mem0_183_4, 
        p_wishbone_bd_ram_mem0_183_5, p_wishbone_bd_ram_mem0_183_6, 
        p_wishbone_bd_ram_mem0_183_7, p_wishbone_bd_ram_mem0_184_0, 
        p_wishbone_bd_ram_mem0_184_1, p_wishbone_bd_ram_mem0_184_2, 
        p_wishbone_bd_ram_mem0_184_3, p_wishbone_bd_ram_mem0_184_4, 
        p_wishbone_bd_ram_mem0_184_5, p_wishbone_bd_ram_mem0_184_6, 
        p_wishbone_bd_ram_mem0_184_7, p_wishbone_bd_ram_mem0_185_0, 
        p_wishbone_bd_ram_mem0_185_1, p_wishbone_bd_ram_mem0_185_2, 
        p_wishbone_bd_ram_mem0_185_3, p_wishbone_bd_ram_mem0_185_4, 
        p_wishbone_bd_ram_mem0_185_5, p_wishbone_bd_ram_mem0_185_6, 
        p_wishbone_bd_ram_mem0_185_7, p_wishbone_bd_ram_mem0_186_0, 
        p_wishbone_bd_ram_mem0_186_1, p_wishbone_bd_ram_mem0_186_2, 
        p_wishbone_bd_ram_mem0_186_3, p_wishbone_bd_ram_mem0_186_4, 
        p_wishbone_bd_ram_mem0_186_5, p_wishbone_bd_ram_mem0_186_6, 
        p_wishbone_bd_ram_mem0_186_7, p_wishbone_bd_ram_mem0_187_0, 
        p_wishbone_bd_ram_mem0_187_1, p_wishbone_bd_ram_mem0_187_2, 
        p_wishbone_bd_ram_mem0_187_3, p_wishbone_bd_ram_mem0_187_4, 
        p_wishbone_bd_ram_mem0_187_5, p_wishbone_bd_ram_mem0_187_6, 
        p_wishbone_bd_ram_mem0_187_7, p_wishbone_bd_ram_mem0_188_0, 
        p_wishbone_bd_ram_mem0_188_1, p_wishbone_bd_ram_mem0_188_2, 
        p_wishbone_bd_ram_mem0_188_3, p_wishbone_bd_ram_mem0_188_4, 
        p_wishbone_bd_ram_mem0_188_5, p_wishbone_bd_ram_mem0_188_6, 
        p_wishbone_bd_ram_mem0_188_7, p_wishbone_bd_ram_mem0_189_0, 
        p_wishbone_bd_ram_mem0_189_1, p_wishbone_bd_ram_mem0_189_2, 
        p_wishbone_bd_ram_mem0_189_3, p_wishbone_bd_ram_mem0_189_4, 
        p_wishbone_bd_ram_mem0_189_5, p_wishbone_bd_ram_mem0_189_6, 
        p_wishbone_bd_ram_mem0_189_7, p_wishbone_bd_ram_mem0_190_0, 
        p_wishbone_bd_ram_mem0_190_1, p_wishbone_bd_ram_mem0_190_2, 
        p_wishbone_bd_ram_mem0_190_3, p_wishbone_bd_ram_mem0_190_4, 
        p_wishbone_bd_ram_mem0_190_5, p_wishbone_bd_ram_mem0_190_6, 
        p_wishbone_bd_ram_mem0_190_7, p_wishbone_bd_ram_mem0_191_0, 
        p_wishbone_bd_ram_mem0_191_1, p_wishbone_bd_ram_mem0_191_2, 
        p_wishbone_bd_ram_mem0_191_3, p_wishbone_bd_ram_mem0_191_4, 
        p_wishbone_bd_ram_mem0_191_5, p_wishbone_bd_ram_mem0_191_6, 
        p_wishbone_bd_ram_mem0_191_7, p_wishbone_bd_ram_mem0_192_0, 
        p_wishbone_bd_ram_mem0_192_1, p_wishbone_bd_ram_mem0_192_2, 
        p_wishbone_bd_ram_mem0_192_3, p_wishbone_bd_ram_mem0_192_4, 
        p_wishbone_bd_ram_mem0_192_5, p_wishbone_bd_ram_mem0_192_6, 
        p_wishbone_bd_ram_mem0_192_7, p_wishbone_bd_ram_mem0_193_0, 
        p_wishbone_bd_ram_mem0_193_1, p_wishbone_bd_ram_mem0_193_2, 
        p_wishbone_bd_ram_mem0_193_3, p_wishbone_bd_ram_mem0_193_4, 
        p_wishbone_bd_ram_mem0_193_5, p_wishbone_bd_ram_mem0_193_6, 
        p_wishbone_bd_ram_mem0_193_7, p_wishbone_bd_ram_mem0_194_0, 
        p_wishbone_bd_ram_mem0_194_1, p_wishbone_bd_ram_mem0_194_2, 
        p_wishbone_bd_ram_mem0_194_3, p_wishbone_bd_ram_mem0_194_4, 
        p_wishbone_bd_ram_mem0_194_5, p_wishbone_bd_ram_mem0_194_6, 
        p_wishbone_bd_ram_mem0_194_7, p_wishbone_bd_ram_mem0_195_0, 
        p_wishbone_bd_ram_mem0_195_1, p_wishbone_bd_ram_mem0_195_2, 
        p_wishbone_bd_ram_mem0_195_3, p_wishbone_bd_ram_mem0_195_4, 
        p_wishbone_bd_ram_mem0_195_5, p_wishbone_bd_ram_mem0_195_6, 
        p_wishbone_bd_ram_mem0_195_7, p_wishbone_bd_ram_mem0_196_0, 
        p_wishbone_bd_ram_mem0_196_1, p_wishbone_bd_ram_mem0_196_2, 
        p_wishbone_bd_ram_mem0_196_3, p_wishbone_bd_ram_mem0_196_4, 
        p_wishbone_bd_ram_mem0_196_5, p_wishbone_bd_ram_mem0_196_6, 
        p_wishbone_bd_ram_mem0_196_7, p_wishbone_bd_ram_mem0_197_0, 
        p_wishbone_bd_ram_mem0_197_1, p_wishbone_bd_ram_mem0_197_2, 
        p_wishbone_bd_ram_mem0_197_3, p_wishbone_bd_ram_mem0_197_4, 
        p_wishbone_bd_ram_mem0_197_5, p_wishbone_bd_ram_mem0_197_6, 
        p_wishbone_bd_ram_mem0_197_7, p_wishbone_bd_ram_mem0_198_0, 
        p_wishbone_bd_ram_mem0_198_1, p_wishbone_bd_ram_mem0_198_2, 
        p_wishbone_bd_ram_mem0_198_3, p_wishbone_bd_ram_mem0_198_4, 
        p_wishbone_bd_ram_mem0_198_5, p_wishbone_bd_ram_mem0_198_6, 
        p_wishbone_bd_ram_mem0_198_7, p_wishbone_bd_ram_mem0_199_0, 
        p_wishbone_bd_ram_mem0_199_1, p_wishbone_bd_ram_mem0_199_2, 
        p_wishbone_bd_ram_mem0_199_3, p_wishbone_bd_ram_mem0_199_4, 
        p_wishbone_bd_ram_mem0_199_5, p_wishbone_bd_ram_mem0_199_6, 
        p_wishbone_bd_ram_mem0_199_7, p_wishbone_bd_ram_mem0_200_0, 
        p_wishbone_bd_ram_mem0_200_1, p_wishbone_bd_ram_mem0_200_2, 
        p_wishbone_bd_ram_mem0_200_3, p_wishbone_bd_ram_mem0_200_4, 
        p_wishbone_bd_ram_mem0_200_5, p_wishbone_bd_ram_mem0_200_6, 
        p_wishbone_bd_ram_mem0_200_7, p_wishbone_bd_ram_mem0_201_0, 
        p_wishbone_bd_ram_mem0_201_1, p_wishbone_bd_ram_mem0_201_2, 
        p_wishbone_bd_ram_mem0_201_3, p_wishbone_bd_ram_mem0_201_4, 
        p_wishbone_bd_ram_mem0_201_5, p_wishbone_bd_ram_mem0_201_6, 
        p_wishbone_bd_ram_mem0_201_7, p_wishbone_bd_ram_mem0_202_0, 
        p_wishbone_bd_ram_mem0_202_1, p_wishbone_bd_ram_mem0_202_2, 
        p_wishbone_bd_ram_mem0_202_3, p_wishbone_bd_ram_mem0_202_4, 
        p_wishbone_bd_ram_mem0_202_5, p_wishbone_bd_ram_mem0_202_6, 
        p_wishbone_bd_ram_mem0_202_7, p_wishbone_bd_ram_mem0_203_0, 
        p_wishbone_bd_ram_mem0_203_1, p_wishbone_bd_ram_mem0_203_2, 
        p_wishbone_bd_ram_mem0_203_3, p_wishbone_bd_ram_mem0_203_4, 
        p_wishbone_bd_ram_mem0_203_5, p_wishbone_bd_ram_mem0_203_6, 
        p_wishbone_bd_ram_mem0_203_7, p_wishbone_bd_ram_mem0_204_0, 
        p_wishbone_bd_ram_mem0_204_1, p_wishbone_bd_ram_mem0_204_2, 
        p_wishbone_bd_ram_mem0_204_3, p_wishbone_bd_ram_mem0_204_4, 
        p_wishbone_bd_ram_mem0_204_5, p_wishbone_bd_ram_mem0_204_6, 
        p_wishbone_bd_ram_mem0_204_7, p_wishbone_bd_ram_mem0_205_0, 
        p_wishbone_bd_ram_mem0_205_1, p_wishbone_bd_ram_mem0_205_2, 
        p_wishbone_bd_ram_mem0_205_3, p_wishbone_bd_ram_mem0_205_4, 
        p_wishbone_bd_ram_mem0_205_5, p_wishbone_bd_ram_mem0_205_6, 
        p_wishbone_bd_ram_mem0_205_7, p_wishbone_bd_ram_mem0_206_0, 
        p_wishbone_bd_ram_mem0_206_1, p_wishbone_bd_ram_mem0_206_2, 
        p_wishbone_bd_ram_mem0_206_3, p_wishbone_bd_ram_mem0_206_4, 
        p_wishbone_bd_ram_mem0_206_5, p_wishbone_bd_ram_mem0_206_6, 
        p_wishbone_bd_ram_mem0_206_7, p_wishbone_bd_ram_mem0_207_0, 
        p_wishbone_bd_ram_mem0_207_1, p_wishbone_bd_ram_mem0_207_2, 
        p_wishbone_bd_ram_mem0_207_3, p_wishbone_bd_ram_mem0_207_4, 
        p_wishbone_bd_ram_mem0_207_5, p_wishbone_bd_ram_mem0_207_6, 
        p_wishbone_bd_ram_mem0_207_7, p_wishbone_bd_ram_mem0_208_0, 
        p_wishbone_bd_ram_mem0_208_1, p_wishbone_bd_ram_mem0_208_2, 
        p_wishbone_bd_ram_mem0_208_3, p_wishbone_bd_ram_mem0_208_4, 
        p_wishbone_bd_ram_mem0_208_5, p_wishbone_bd_ram_mem0_208_6, 
        p_wishbone_bd_ram_mem0_208_7, p_wishbone_bd_ram_mem0_209_0, 
        p_wishbone_bd_ram_mem0_209_1, p_wishbone_bd_ram_mem0_209_2, 
        p_wishbone_bd_ram_mem0_209_3, p_wishbone_bd_ram_mem0_209_4, 
        p_wishbone_bd_ram_mem0_209_5, p_wishbone_bd_ram_mem0_209_6, 
        p_wishbone_bd_ram_mem0_209_7, p_wishbone_bd_ram_mem0_210_0, 
        p_wishbone_bd_ram_mem0_210_1, p_wishbone_bd_ram_mem0_210_2, 
        p_wishbone_bd_ram_mem0_210_3, p_wishbone_bd_ram_mem0_210_4, 
        p_wishbone_bd_ram_mem0_210_5, p_wishbone_bd_ram_mem0_210_6, 
        p_wishbone_bd_ram_mem0_210_7, p_wishbone_bd_ram_mem0_211_0, 
        p_wishbone_bd_ram_mem0_211_1, p_wishbone_bd_ram_mem0_211_2, 
        p_wishbone_bd_ram_mem0_211_3, p_wishbone_bd_ram_mem0_211_4, 
        p_wishbone_bd_ram_mem0_211_5, p_wishbone_bd_ram_mem0_211_6, 
        p_wishbone_bd_ram_mem0_211_7, p_wishbone_bd_ram_mem0_212_0, 
        p_wishbone_bd_ram_mem0_212_1, p_wishbone_bd_ram_mem0_212_2, 
        p_wishbone_bd_ram_mem0_212_3, p_wishbone_bd_ram_mem0_212_4, 
        p_wishbone_bd_ram_mem0_212_5, p_wishbone_bd_ram_mem0_212_6, 
        p_wishbone_bd_ram_mem0_212_7, p_wishbone_bd_ram_mem0_213_0, 
        p_wishbone_bd_ram_mem0_213_1, p_wishbone_bd_ram_mem0_213_2, 
        p_wishbone_bd_ram_mem0_213_3, p_wishbone_bd_ram_mem0_213_4, 
        p_wishbone_bd_ram_mem0_213_5, p_wishbone_bd_ram_mem0_213_6, 
        p_wishbone_bd_ram_mem0_213_7, p_wishbone_bd_ram_mem0_214_0, 
        p_wishbone_bd_ram_mem0_214_1, p_wishbone_bd_ram_mem0_214_2, 
        p_wishbone_bd_ram_mem0_214_3, p_wishbone_bd_ram_mem0_214_4, 
        p_wishbone_bd_ram_mem0_214_5, p_wishbone_bd_ram_mem0_214_6, 
        p_wishbone_bd_ram_mem0_214_7, p_wishbone_bd_ram_mem0_215_0, 
        p_wishbone_bd_ram_mem0_215_1, p_wishbone_bd_ram_mem0_215_2, 
        p_wishbone_bd_ram_mem0_215_3, p_wishbone_bd_ram_mem0_215_4, 
        p_wishbone_bd_ram_mem0_215_5, p_wishbone_bd_ram_mem0_215_6, 
        p_wishbone_bd_ram_mem0_215_7, p_wishbone_bd_ram_mem0_216_0, 
        p_wishbone_bd_ram_mem0_216_1, p_wishbone_bd_ram_mem0_216_2, 
        p_wishbone_bd_ram_mem0_216_3, p_wishbone_bd_ram_mem0_216_4, 
        p_wishbone_bd_ram_mem0_216_5, p_wishbone_bd_ram_mem0_216_6, 
        p_wishbone_bd_ram_mem0_216_7, p_wishbone_bd_ram_mem0_217_0, 
        p_wishbone_bd_ram_mem0_217_1, p_wishbone_bd_ram_mem0_217_2, 
        p_wishbone_bd_ram_mem0_217_3, p_wishbone_bd_ram_mem0_217_4, 
        p_wishbone_bd_ram_mem0_217_5, p_wishbone_bd_ram_mem0_217_6, 
        p_wishbone_bd_ram_mem0_217_7, p_wishbone_bd_ram_mem0_218_0, 
        p_wishbone_bd_ram_mem0_218_1, p_wishbone_bd_ram_mem0_218_2, 
        p_wishbone_bd_ram_mem0_218_3, p_wishbone_bd_ram_mem0_218_4, 
        p_wishbone_bd_ram_mem0_218_5, p_wishbone_bd_ram_mem0_218_6, 
        p_wishbone_bd_ram_mem0_218_7, p_wishbone_bd_ram_mem0_219_0, 
        p_wishbone_bd_ram_mem0_219_1, p_wishbone_bd_ram_mem0_219_2, 
        p_wishbone_bd_ram_mem0_219_3, p_wishbone_bd_ram_mem0_219_4, 
        p_wishbone_bd_ram_mem0_219_5, p_wishbone_bd_ram_mem0_219_6, 
        p_wishbone_bd_ram_mem0_219_7, p_wishbone_bd_ram_mem0_220_0, 
        p_wishbone_bd_ram_mem0_220_1, p_wishbone_bd_ram_mem0_220_2, 
        p_wishbone_bd_ram_mem0_220_3, p_wishbone_bd_ram_mem0_220_4, 
        p_wishbone_bd_ram_mem0_220_5, p_wishbone_bd_ram_mem0_220_6, 
        p_wishbone_bd_ram_mem0_220_7, p_wishbone_bd_ram_mem0_221_0, 
        p_wishbone_bd_ram_mem0_221_1, p_wishbone_bd_ram_mem0_221_2, 
        p_wishbone_bd_ram_mem0_221_3, p_wishbone_bd_ram_mem0_221_4, 
        p_wishbone_bd_ram_mem0_221_5, p_wishbone_bd_ram_mem0_221_6, 
        p_wishbone_bd_ram_mem0_221_7, p_wishbone_bd_ram_mem0_222_0, 
        p_wishbone_bd_ram_mem0_222_1, p_wishbone_bd_ram_mem0_222_2, 
        p_wishbone_bd_ram_mem0_222_3, p_wishbone_bd_ram_mem0_222_4, 
        p_wishbone_bd_ram_mem0_222_5, p_wishbone_bd_ram_mem0_222_6, 
        p_wishbone_bd_ram_mem0_222_7, p_wishbone_bd_ram_mem0_223_0, 
        p_wishbone_bd_ram_mem0_223_1, p_wishbone_bd_ram_mem0_223_2, 
        p_wishbone_bd_ram_mem0_223_3, p_wishbone_bd_ram_mem0_223_4, 
        p_wishbone_bd_ram_mem0_223_5, p_wishbone_bd_ram_mem0_223_6, 
        p_wishbone_bd_ram_mem0_223_7, p_wishbone_bd_ram_mem0_224_0, 
        p_wishbone_bd_ram_mem0_224_1, p_wishbone_bd_ram_mem0_224_2, 
        p_wishbone_bd_ram_mem0_224_3, p_wishbone_bd_ram_mem0_224_4, 
        p_wishbone_bd_ram_mem0_224_5, p_wishbone_bd_ram_mem0_224_6, 
        p_wishbone_bd_ram_mem0_224_7, p_wishbone_bd_ram_mem0_225_0, 
        p_wishbone_bd_ram_mem0_225_1, p_wishbone_bd_ram_mem0_225_2, 
        p_wishbone_bd_ram_mem0_225_3, p_wishbone_bd_ram_mem0_225_4, 
        p_wishbone_bd_ram_mem0_225_5, p_wishbone_bd_ram_mem0_225_6, 
        p_wishbone_bd_ram_mem0_225_7, p_wishbone_bd_ram_mem0_226_0, 
        p_wishbone_bd_ram_mem0_226_1, p_wishbone_bd_ram_mem0_226_2, 
        p_wishbone_bd_ram_mem0_226_3, p_wishbone_bd_ram_mem0_226_4, 
        p_wishbone_bd_ram_mem0_226_5, p_wishbone_bd_ram_mem0_226_6, 
        p_wishbone_bd_ram_mem0_226_7, p_wishbone_bd_ram_mem0_227_0, 
        p_wishbone_bd_ram_mem0_227_1, p_wishbone_bd_ram_mem0_227_2, 
        p_wishbone_bd_ram_mem0_227_3, p_wishbone_bd_ram_mem0_227_4, 
        p_wishbone_bd_ram_mem0_227_5, p_wishbone_bd_ram_mem0_227_6, 
        p_wishbone_bd_ram_mem0_227_7, p_wishbone_bd_ram_mem0_228_0, 
        p_wishbone_bd_ram_mem0_228_1, p_wishbone_bd_ram_mem0_228_2, 
        p_wishbone_bd_ram_mem0_228_3, p_wishbone_bd_ram_mem0_228_4, 
        p_wishbone_bd_ram_mem0_228_5, p_wishbone_bd_ram_mem0_228_6, 
        p_wishbone_bd_ram_mem0_228_7, p_wishbone_bd_ram_mem0_229_0, 
        p_wishbone_bd_ram_mem0_229_1, p_wishbone_bd_ram_mem0_229_2, 
        p_wishbone_bd_ram_mem0_229_3, p_wishbone_bd_ram_mem0_229_4, 
        p_wishbone_bd_ram_mem0_229_5, p_wishbone_bd_ram_mem0_229_6, 
        p_wishbone_bd_ram_mem0_229_7, p_wishbone_bd_ram_mem0_230_0, 
        p_wishbone_bd_ram_mem0_230_1, p_wishbone_bd_ram_mem0_230_2, 
        p_wishbone_bd_ram_mem0_230_3, p_wishbone_bd_ram_mem0_230_4, 
        p_wishbone_bd_ram_mem0_230_5, p_wishbone_bd_ram_mem0_230_6, 
        p_wishbone_bd_ram_mem0_230_7, p_wishbone_bd_ram_mem0_231_0, 
        p_wishbone_bd_ram_mem0_231_1, p_wishbone_bd_ram_mem0_231_2, 
        p_wishbone_bd_ram_mem0_231_3, p_wishbone_bd_ram_mem0_231_4, 
        p_wishbone_bd_ram_mem0_231_5, p_wishbone_bd_ram_mem0_231_6, 
        p_wishbone_bd_ram_mem0_231_7, p_wishbone_bd_ram_mem0_232_0, 
        p_wishbone_bd_ram_mem0_232_1, p_wishbone_bd_ram_mem0_232_2, 
        p_wishbone_bd_ram_mem0_232_3, p_wishbone_bd_ram_mem0_232_4, 
        p_wishbone_bd_ram_mem0_232_5, p_wishbone_bd_ram_mem0_232_6, 
        p_wishbone_bd_ram_mem0_232_7, p_wishbone_bd_ram_mem0_233_0, 
        p_wishbone_bd_ram_mem0_233_1, p_wishbone_bd_ram_mem0_233_2, 
        p_wishbone_bd_ram_mem0_233_3, p_wishbone_bd_ram_mem0_233_4, 
        p_wishbone_bd_ram_mem0_233_5, p_wishbone_bd_ram_mem0_233_6, 
        p_wishbone_bd_ram_mem0_233_7, p_wishbone_bd_ram_mem0_234_0, 
        p_wishbone_bd_ram_mem0_234_1, p_wishbone_bd_ram_mem0_234_2, 
        p_wishbone_bd_ram_mem0_234_3, p_wishbone_bd_ram_mem0_234_4, 
        p_wishbone_bd_ram_mem0_234_5, p_wishbone_bd_ram_mem0_234_6, 
        p_wishbone_bd_ram_mem0_234_7, p_wishbone_bd_ram_mem0_235_0, 
        p_wishbone_bd_ram_mem0_235_1, p_wishbone_bd_ram_mem0_235_2, 
        p_wishbone_bd_ram_mem0_235_3, p_wishbone_bd_ram_mem0_235_4, 
        p_wishbone_bd_ram_mem0_235_5, p_wishbone_bd_ram_mem0_235_6, 
        p_wishbone_bd_ram_mem0_235_7, p_wishbone_bd_ram_mem0_236_0, 
        p_wishbone_bd_ram_mem0_236_1, p_wishbone_bd_ram_mem0_236_2, 
        p_wishbone_bd_ram_mem0_236_3, p_wishbone_bd_ram_mem0_236_4, 
        p_wishbone_bd_ram_mem0_236_5, p_wishbone_bd_ram_mem0_236_6, 
        p_wishbone_bd_ram_mem0_236_7, p_wishbone_bd_ram_mem0_237_0, 
        p_wishbone_bd_ram_mem0_237_1, p_wishbone_bd_ram_mem0_237_2, 
        p_wishbone_bd_ram_mem0_237_3, p_wishbone_bd_ram_mem0_237_4, 
        p_wishbone_bd_ram_mem0_237_5, p_wishbone_bd_ram_mem0_237_6, 
        p_wishbone_bd_ram_mem0_237_7, p_wishbone_bd_ram_mem0_238_0, 
        p_wishbone_bd_ram_mem0_238_1, p_wishbone_bd_ram_mem0_238_2, 
        p_wishbone_bd_ram_mem0_238_3, p_wishbone_bd_ram_mem0_238_4, 
        p_wishbone_bd_ram_mem0_238_5, p_wishbone_bd_ram_mem0_238_6, 
        p_wishbone_bd_ram_mem0_238_7, p_wishbone_bd_ram_mem0_239_0, 
        p_wishbone_bd_ram_mem0_239_1, p_wishbone_bd_ram_mem0_239_2, 
        p_wishbone_bd_ram_mem0_239_3, p_wishbone_bd_ram_mem0_239_4, 
        p_wishbone_bd_ram_mem0_239_5, p_wishbone_bd_ram_mem0_239_6, 
        p_wishbone_bd_ram_mem0_239_7, p_wishbone_bd_ram_mem0_240_0, 
        p_wishbone_bd_ram_mem0_240_1, p_wishbone_bd_ram_mem0_240_2, 
        p_wishbone_bd_ram_mem0_240_3, p_wishbone_bd_ram_mem0_240_4, 
        p_wishbone_bd_ram_mem0_240_5, p_wishbone_bd_ram_mem0_240_6, 
        p_wishbone_bd_ram_mem0_240_7, p_wishbone_bd_ram_mem0_241_0, 
        p_wishbone_bd_ram_mem0_241_1, p_wishbone_bd_ram_mem0_241_2, 
        p_wishbone_bd_ram_mem0_241_3, p_wishbone_bd_ram_mem0_241_4, 
        p_wishbone_bd_ram_mem0_241_5, p_wishbone_bd_ram_mem0_241_6, 
        p_wishbone_bd_ram_mem0_241_7, p_wishbone_bd_ram_mem0_242_0, 
        p_wishbone_bd_ram_mem0_242_1, p_wishbone_bd_ram_mem0_242_2, 
        p_wishbone_bd_ram_mem0_242_3, p_wishbone_bd_ram_mem0_242_4, 
        p_wishbone_bd_ram_mem0_242_5, p_wishbone_bd_ram_mem0_242_6, 
        p_wishbone_bd_ram_mem0_242_7, p_wishbone_bd_ram_mem0_243_0, 
        p_wishbone_bd_ram_mem0_243_1, p_wishbone_bd_ram_mem0_243_2, 
        p_wishbone_bd_ram_mem0_243_3, p_wishbone_bd_ram_mem0_243_4, 
        p_wishbone_bd_ram_mem0_243_5, p_wishbone_bd_ram_mem0_243_6, 
        p_wishbone_bd_ram_mem0_243_7, p_wishbone_bd_ram_mem0_244_0, 
        p_wishbone_bd_ram_mem0_244_1, p_wishbone_bd_ram_mem0_244_2, 
        p_wishbone_bd_ram_mem0_244_3, p_wishbone_bd_ram_mem0_244_4, 
        p_wishbone_bd_ram_mem0_244_5, p_wishbone_bd_ram_mem0_244_6, 
        p_wishbone_bd_ram_mem0_244_7, p_wishbone_bd_ram_mem0_245_0, 
        p_wishbone_bd_ram_mem0_245_1, p_wishbone_bd_ram_mem0_245_2, 
        p_wishbone_bd_ram_mem0_245_3, p_wishbone_bd_ram_mem0_245_4, 
        p_wishbone_bd_ram_mem0_245_5, p_wishbone_bd_ram_mem0_245_6, 
        p_wishbone_bd_ram_mem0_245_7, p_wishbone_bd_ram_mem0_246_0, 
        p_wishbone_bd_ram_mem0_246_1, p_wishbone_bd_ram_mem0_246_2, 
        p_wishbone_bd_ram_mem0_246_3, p_wishbone_bd_ram_mem0_246_4, 
        p_wishbone_bd_ram_mem0_246_5, p_wishbone_bd_ram_mem0_246_6, 
        p_wishbone_bd_ram_mem0_246_7, p_wishbone_bd_ram_mem0_247_0, 
        p_wishbone_bd_ram_mem0_247_1, p_wishbone_bd_ram_mem0_247_2, 
        p_wishbone_bd_ram_mem0_247_3, p_wishbone_bd_ram_mem0_247_4, 
        p_wishbone_bd_ram_mem0_247_5, p_wishbone_bd_ram_mem0_247_6, 
        p_wishbone_bd_ram_mem0_247_7, p_wishbone_bd_ram_mem0_248_0, 
        p_wishbone_bd_ram_mem0_248_1, p_wishbone_bd_ram_mem0_248_2, 
        p_wishbone_bd_ram_mem0_248_3, p_wishbone_bd_ram_mem0_248_4, 
        p_wishbone_bd_ram_mem0_248_5, p_wishbone_bd_ram_mem0_248_6, 
        p_wishbone_bd_ram_mem0_248_7, p_wishbone_bd_ram_mem0_249_0, 
        p_wishbone_bd_ram_mem0_249_1, p_wishbone_bd_ram_mem0_249_2, 
        p_wishbone_bd_ram_mem0_249_3, p_wishbone_bd_ram_mem0_249_4, 
        p_wishbone_bd_ram_mem0_249_5, p_wishbone_bd_ram_mem0_249_6, 
        p_wishbone_bd_ram_mem0_249_7, p_wishbone_bd_ram_mem0_250_0, 
        p_wishbone_bd_ram_mem0_250_1, p_wishbone_bd_ram_mem0_250_2, 
        p_wishbone_bd_ram_mem0_250_3, p_wishbone_bd_ram_mem0_250_4, 
        p_wishbone_bd_ram_mem0_250_5, p_wishbone_bd_ram_mem0_250_6, 
        p_wishbone_bd_ram_mem0_250_7, p_wishbone_bd_ram_mem0_251_0, 
        p_wishbone_bd_ram_mem0_251_1, p_wishbone_bd_ram_mem0_251_2, 
        p_wishbone_bd_ram_mem0_251_3, p_wishbone_bd_ram_mem0_251_4, 
        p_wishbone_bd_ram_mem0_251_5, p_wishbone_bd_ram_mem0_251_6, 
        p_wishbone_bd_ram_mem0_251_7, p_wishbone_bd_ram_mem0_252_0, 
        p_wishbone_bd_ram_mem0_252_1, p_wishbone_bd_ram_mem0_252_2, 
        p_wishbone_bd_ram_mem0_252_3, p_wishbone_bd_ram_mem0_252_4, 
        p_wishbone_bd_ram_mem0_252_5, p_wishbone_bd_ram_mem0_252_6, 
        p_wishbone_bd_ram_mem0_252_7, p_wishbone_bd_ram_mem0_253_0, 
        p_wishbone_bd_ram_mem0_253_1, p_wishbone_bd_ram_mem0_253_2, 
        p_wishbone_bd_ram_mem0_253_3, p_wishbone_bd_ram_mem0_253_4, 
        p_wishbone_bd_ram_mem0_253_5, p_wishbone_bd_ram_mem0_253_6, 
        p_wishbone_bd_ram_mem0_253_7, p_wishbone_bd_ram_mem0_254_0, 
        p_wishbone_bd_ram_mem0_254_1, p_wishbone_bd_ram_mem0_254_2, 
        p_wishbone_bd_ram_mem0_254_3, p_wishbone_bd_ram_mem0_254_4, 
        p_wishbone_bd_ram_mem0_254_5, p_wishbone_bd_ram_mem0_254_6, 
        p_wishbone_bd_ram_mem0_254_7, p_wishbone_bd_ram_mem0_255_0, 
        p_wishbone_bd_ram_mem0_255_1, p_wishbone_bd_ram_mem0_255_2, 
        p_wishbone_bd_ram_mem0_255_3, p_wishbone_bd_ram_mem0_255_4, 
        p_wishbone_bd_ram_mem0_255_5, p_wishbone_bd_ram_mem0_255_6, 
        p_wishbone_bd_ram_mem0_255_7, p_wishbone_bd_ram_N102, 
        p_wishbone_bd_ram_N103, p_wishbone_bd_ram_N104, p_wishbone_bd_ram_N105, 
        p_wishbone_bd_ram_N106, p_wishbone_bd_ram_N107, p_wishbone_bd_ram_N108, 
        p_wishbone_bd_ram_N109, p_wishbone_TxData_wb_0, p_wishbone_TxData_wb_1, 
        p_wishbone_TxData_wb_2, p_wishbone_TxData_wb_3, p_wishbone_TxData_wb_4, 
        p_wishbone_TxData_wb_5, p_wishbone_TxData_wb_6, p_wishbone_TxData_wb_7, 
        p_wishbone_TxData_wb_8, p_wishbone_TxData_wb_9, 
        p_wishbone_TxData_wb_10, p_wishbone_TxData_wb_11, 
        p_wishbone_TxData_wb_12, p_wishbone_TxData_wb_13, 
        p_wishbone_TxData_wb_14, p_wishbone_TxData_wb_15, 
        p_wishbone_TxData_wb_16, p_wishbone_TxData_wb_17, 
        p_wishbone_TxData_wb_18, p_wishbone_TxData_wb_19, 
        p_wishbone_TxData_wb_20, p_wishbone_TxData_wb_21, 
        p_wishbone_TxData_wb_22, p_wishbone_TxData_wb_23, 
        p_wishbone_TxData_wb_24, p_wishbone_TxData_wb_25, 
        p_wishbone_TxData_wb_26, p_wishbone_TxData_wb_27, 
        p_wishbone_TxData_wb_28, p_wishbone_TxData_wb_29, 
        p_wishbone_TxData_wb_30, p_wishbone_TxData_wb_31, 
        p_wishbone_tx_fifo_fifo_15_0, p_wishbone_tx_fifo_fifo_15_1, 
        p_wishbone_tx_fifo_fifo_15_2, p_wishbone_tx_fifo_fifo_15_3, 
        p_wishbone_tx_fifo_fifo_15_4, p_wishbone_tx_fifo_fifo_15_5, 
        p_wishbone_tx_fifo_fifo_15_6, p_wishbone_tx_fifo_fifo_15_7, 
        p_wishbone_tx_fifo_fifo_15_8, p_wishbone_tx_fifo_fifo_15_9, 
        p_wishbone_tx_fifo_fifo_15_10, p_wishbone_tx_fifo_fifo_15_11, 
        p_wishbone_tx_fifo_fifo_15_12, p_wishbone_tx_fifo_fifo_15_13, 
        p_wishbone_tx_fifo_fifo_15_14, p_wishbone_tx_fifo_fifo_15_15, 
        p_wishbone_tx_fifo_fifo_15_16, p_wishbone_tx_fifo_fifo_15_17, 
        p_wishbone_tx_fifo_fifo_15_18, p_wishbone_tx_fifo_fifo_15_19, 
        p_wishbone_tx_fifo_fifo_15_20, p_wishbone_tx_fifo_fifo_15_21, 
        p_wishbone_tx_fifo_fifo_15_22, p_wishbone_tx_fifo_fifo_15_23, 
        p_wishbone_tx_fifo_fifo_15_24, p_wishbone_tx_fifo_fifo_15_25, 
        p_wishbone_tx_fifo_fifo_15_26, p_wishbone_tx_fifo_fifo_15_27, 
        p_wishbone_tx_fifo_fifo_15_28, p_wishbone_tx_fifo_fifo_15_29, 
        p_wishbone_tx_fifo_fifo_15_30, p_wishbone_tx_fifo_fifo_15_31, 
        p_wishbone_tx_fifo_fifo_14_0, p_wishbone_tx_fifo_fifo_14_1, 
        p_wishbone_tx_fifo_fifo_14_2, p_wishbone_tx_fifo_fifo_14_3, 
        p_wishbone_tx_fifo_fifo_14_4, p_wishbone_tx_fifo_fifo_14_5, 
        p_wishbone_tx_fifo_fifo_14_6, p_wishbone_tx_fifo_fifo_14_7, 
        p_wishbone_tx_fifo_fifo_14_8, p_wishbone_tx_fifo_fifo_14_9, 
        p_wishbone_tx_fifo_fifo_14_10, p_wishbone_tx_fifo_fifo_14_11, 
        p_wishbone_tx_fifo_fifo_14_12, p_wishbone_tx_fifo_fifo_14_13, 
        p_wishbone_tx_fifo_fifo_14_14, p_wishbone_tx_fifo_fifo_14_15, 
        p_wishbone_tx_fifo_fifo_14_16, p_wishbone_tx_fifo_fifo_14_17, 
        p_wishbone_tx_fifo_fifo_14_18, p_wishbone_tx_fifo_fifo_14_19, 
        p_wishbone_tx_fifo_fifo_14_20, p_wishbone_tx_fifo_fifo_14_21, 
        p_wishbone_tx_fifo_fifo_14_22, p_wishbone_tx_fifo_fifo_14_23, 
        p_wishbone_tx_fifo_fifo_14_24, p_wishbone_tx_fifo_fifo_14_25, 
        p_wishbone_tx_fifo_fifo_14_26, p_wishbone_tx_fifo_fifo_14_27, 
        p_wishbone_tx_fifo_fifo_14_28, p_wishbone_tx_fifo_fifo_14_29, 
        p_wishbone_tx_fifo_fifo_14_30, p_wishbone_tx_fifo_fifo_14_31, 
        p_wishbone_tx_fifo_fifo_13_0, p_wishbone_tx_fifo_fifo_13_1, 
        p_wishbone_tx_fifo_fifo_13_2, p_wishbone_tx_fifo_fifo_13_3, 
        p_wishbone_tx_fifo_fifo_13_4, p_wishbone_tx_fifo_fifo_13_5, 
        p_wishbone_tx_fifo_fifo_13_6, p_wishbone_tx_fifo_fifo_13_7, 
        p_wishbone_tx_fifo_fifo_13_8, p_wishbone_tx_fifo_fifo_13_9, 
        p_wishbone_tx_fifo_fifo_13_10, p_wishbone_tx_fifo_fifo_13_11, 
        p_wishbone_tx_fifo_fifo_13_12, p_wishbone_tx_fifo_fifo_13_13, 
        p_wishbone_tx_fifo_fifo_13_14, p_wishbone_tx_fifo_fifo_13_15, 
        p_wishbone_tx_fifo_fifo_13_16, p_wishbone_tx_fifo_fifo_13_17, 
        p_wishbone_tx_fifo_fifo_13_18, p_wishbone_tx_fifo_fifo_13_19, 
        p_wishbone_tx_fifo_fifo_13_20, p_wishbone_tx_fifo_fifo_13_21, 
        p_wishbone_tx_fifo_fifo_13_22, p_wishbone_tx_fifo_fifo_13_23, 
        p_wishbone_tx_fifo_fifo_13_24, p_wishbone_tx_fifo_fifo_13_25, 
        p_wishbone_tx_fifo_fifo_13_26, p_wishbone_tx_fifo_fifo_13_27, 
        p_wishbone_tx_fifo_fifo_13_28, p_wishbone_tx_fifo_fifo_13_29, 
        p_wishbone_tx_fifo_fifo_13_30, p_wishbone_tx_fifo_fifo_13_31, 
        p_wishbone_tx_fifo_fifo_12_0, p_wishbone_tx_fifo_fifo_12_1, 
        p_wishbone_tx_fifo_fifo_12_2, p_wishbone_tx_fifo_fifo_12_3, 
        p_wishbone_tx_fifo_fifo_12_4, p_wishbone_tx_fifo_fifo_12_5, 
        p_wishbone_tx_fifo_fifo_12_6, p_wishbone_tx_fifo_fifo_12_7, 
        p_wishbone_tx_fifo_fifo_12_8, p_wishbone_tx_fifo_fifo_12_9, 
        p_wishbone_tx_fifo_fifo_12_10, p_wishbone_tx_fifo_fifo_12_11, 
        p_wishbone_tx_fifo_fifo_12_12, p_wishbone_tx_fifo_fifo_12_13, 
        p_wishbone_tx_fifo_fifo_12_14, p_wishbone_tx_fifo_fifo_12_15, 
        p_wishbone_tx_fifo_fifo_12_16, p_wishbone_tx_fifo_fifo_12_17, 
        p_wishbone_tx_fifo_fifo_12_18, p_wishbone_tx_fifo_fifo_12_19, 
        p_wishbone_tx_fifo_fifo_12_20, p_wishbone_tx_fifo_fifo_12_21, 
        p_wishbone_tx_fifo_fifo_12_22, p_wishbone_tx_fifo_fifo_12_23, 
        p_wishbone_tx_fifo_fifo_12_24, p_wishbone_tx_fifo_fifo_12_25, 
        p_wishbone_tx_fifo_fifo_12_26, p_wishbone_tx_fifo_fifo_12_27, 
        p_wishbone_tx_fifo_fifo_12_28, p_wishbone_tx_fifo_fifo_12_29, 
        p_wishbone_tx_fifo_fifo_12_30, p_wishbone_tx_fifo_fifo_12_31, 
        p_wishbone_tx_fifo_fifo_11_0, p_wishbone_tx_fifo_fifo_11_1, 
        p_wishbone_tx_fifo_fifo_11_2, p_wishbone_tx_fifo_fifo_11_3, 
        p_wishbone_tx_fifo_fifo_11_4, p_wishbone_tx_fifo_fifo_11_5, 
        p_wishbone_tx_fifo_fifo_11_6, p_wishbone_tx_fifo_fifo_11_7, 
        p_wishbone_tx_fifo_fifo_11_8, p_wishbone_tx_fifo_fifo_11_9, 
        p_wishbone_tx_fifo_fifo_11_10, p_wishbone_tx_fifo_fifo_11_11, 
        p_wishbone_tx_fifo_fifo_11_12, p_wishbone_tx_fifo_fifo_11_13, 
        p_wishbone_tx_fifo_fifo_11_14, p_wishbone_tx_fifo_fifo_11_15, 
        p_wishbone_tx_fifo_fifo_11_16, p_wishbone_tx_fifo_fifo_11_17, 
        p_wishbone_tx_fifo_fifo_11_18, p_wishbone_tx_fifo_fifo_11_19, 
        p_wishbone_tx_fifo_fifo_11_20, p_wishbone_tx_fifo_fifo_11_21, 
        p_wishbone_tx_fifo_fifo_11_22, p_wishbone_tx_fifo_fifo_11_23, 
        p_wishbone_tx_fifo_fifo_11_24, p_wishbone_tx_fifo_fifo_11_25, 
        p_wishbone_tx_fifo_fifo_11_26, p_wishbone_tx_fifo_fifo_11_27, 
        p_wishbone_tx_fifo_fifo_11_28, p_wishbone_tx_fifo_fifo_11_29, 
        p_wishbone_tx_fifo_fifo_11_30, p_wishbone_tx_fifo_fifo_11_31, 
        p_wishbone_tx_fifo_fifo_10_0, p_wishbone_tx_fifo_fifo_10_1, 
        p_wishbone_tx_fifo_fifo_10_2, p_wishbone_tx_fifo_fifo_10_3, 
        p_wishbone_tx_fifo_fifo_10_4, p_wishbone_tx_fifo_fifo_10_5, 
        p_wishbone_tx_fifo_fifo_10_6, p_wishbone_tx_fifo_fifo_10_7, 
        p_wishbone_tx_fifo_fifo_10_8, p_wishbone_tx_fifo_fifo_10_9, 
        p_wishbone_tx_fifo_fifo_10_10, p_wishbone_tx_fifo_fifo_10_11, 
        p_wishbone_tx_fifo_fifo_10_12, p_wishbone_tx_fifo_fifo_10_13, 
        p_wishbone_tx_fifo_fifo_10_14, p_wishbone_tx_fifo_fifo_10_15, 
        p_wishbone_tx_fifo_fifo_10_16, p_wishbone_tx_fifo_fifo_10_17, 
        p_wishbone_tx_fifo_fifo_10_18, p_wishbone_tx_fifo_fifo_10_19, 
        p_wishbone_tx_fifo_fifo_10_20, p_wishbone_tx_fifo_fifo_10_21, 
        p_wishbone_tx_fifo_fifo_10_22, p_wishbone_tx_fifo_fifo_10_23, 
        p_wishbone_tx_fifo_fifo_10_24, p_wishbone_tx_fifo_fifo_10_25, 
        p_wishbone_tx_fifo_fifo_10_26, p_wishbone_tx_fifo_fifo_10_27, 
        p_wishbone_tx_fifo_fifo_10_28, p_wishbone_tx_fifo_fifo_10_29, 
        p_wishbone_tx_fifo_fifo_10_30, p_wishbone_tx_fifo_fifo_10_31, 
        p_wishbone_tx_fifo_fifo_9_0, p_wishbone_tx_fifo_fifo_9_1, 
        p_wishbone_tx_fifo_fifo_9_2, p_wishbone_tx_fifo_fifo_9_3, 
        p_wishbone_tx_fifo_fifo_9_4, p_wishbone_tx_fifo_fifo_9_5, 
        p_wishbone_tx_fifo_fifo_9_6, p_wishbone_tx_fifo_fifo_9_7, 
        p_wishbone_tx_fifo_fifo_9_8, p_wishbone_tx_fifo_fifo_9_9, 
        p_wishbone_tx_fifo_fifo_9_10, p_wishbone_tx_fifo_fifo_9_11, 
        p_wishbone_tx_fifo_fifo_9_12, p_wishbone_tx_fifo_fifo_9_13, 
        p_wishbone_tx_fifo_fifo_9_14, p_wishbone_tx_fifo_fifo_9_15, 
        p_wishbone_tx_fifo_fifo_9_16, p_wishbone_tx_fifo_fifo_9_17, 
        p_wishbone_tx_fifo_fifo_9_18, p_wishbone_tx_fifo_fifo_9_19, 
        p_wishbone_tx_fifo_fifo_9_20, p_wishbone_tx_fifo_fifo_9_21, 
        p_wishbone_tx_fifo_fifo_9_22, p_wishbone_tx_fifo_fifo_9_23, 
        p_wishbone_tx_fifo_fifo_9_24, p_wishbone_tx_fifo_fifo_9_25, 
        p_wishbone_tx_fifo_fifo_9_26, p_wishbone_tx_fifo_fifo_9_27, 
        p_wishbone_tx_fifo_fifo_9_28, p_wishbone_tx_fifo_fifo_9_29, 
        p_wishbone_tx_fifo_fifo_9_30, p_wishbone_tx_fifo_fifo_9_31, 
        p_wishbone_tx_fifo_fifo_8_0, p_wishbone_tx_fifo_fifo_8_1, 
        p_wishbone_tx_fifo_fifo_8_2, p_wishbone_tx_fifo_fifo_8_3, 
        p_wishbone_tx_fifo_fifo_8_4, p_wishbone_tx_fifo_fifo_8_5, 
        p_wishbone_tx_fifo_fifo_8_6, p_wishbone_tx_fifo_fifo_8_7, 
        p_wishbone_tx_fifo_fifo_8_8, p_wishbone_tx_fifo_fifo_8_9, 
        p_wishbone_tx_fifo_fifo_8_10, p_wishbone_tx_fifo_fifo_8_11, 
        p_wishbone_tx_fifo_fifo_8_12, p_wishbone_tx_fifo_fifo_8_13, 
        p_wishbone_tx_fifo_fifo_8_14, p_wishbone_tx_fifo_fifo_8_15, 
        p_wishbone_tx_fifo_fifo_8_16, p_wishbone_tx_fifo_fifo_8_17, 
        p_wishbone_tx_fifo_fifo_8_18, p_wishbone_tx_fifo_fifo_8_19, 
        p_wishbone_tx_fifo_fifo_8_20, p_wishbone_tx_fifo_fifo_8_21, 
        p_wishbone_tx_fifo_fifo_8_22, p_wishbone_tx_fifo_fifo_8_23, 
        p_wishbone_tx_fifo_fifo_8_24, p_wishbone_tx_fifo_fifo_8_25, 
        p_wishbone_tx_fifo_fifo_8_26, p_wishbone_tx_fifo_fifo_8_27, 
        p_wishbone_tx_fifo_fifo_8_28, p_wishbone_tx_fifo_fifo_8_29, 
        p_wishbone_tx_fifo_fifo_8_30, p_wishbone_tx_fifo_fifo_8_31, 
        p_wishbone_tx_fifo_fifo_7_0, p_wishbone_tx_fifo_fifo_7_1, 
        p_wishbone_tx_fifo_fifo_7_2, p_wishbone_tx_fifo_fifo_7_3, 
        p_wishbone_tx_fifo_fifo_7_4, p_wishbone_tx_fifo_fifo_7_5, 
        p_wishbone_tx_fifo_fifo_7_6, p_wishbone_tx_fifo_fifo_7_7, 
        p_wishbone_tx_fifo_fifo_7_8, p_wishbone_tx_fifo_fifo_7_9, 
        p_wishbone_tx_fifo_fifo_7_10, p_wishbone_tx_fifo_fifo_7_11, 
        p_wishbone_tx_fifo_fifo_7_12, p_wishbone_tx_fifo_fifo_7_13, 
        p_wishbone_tx_fifo_fifo_7_14, p_wishbone_tx_fifo_fifo_7_15, 
        p_wishbone_tx_fifo_fifo_7_16, p_wishbone_tx_fifo_fifo_7_17, 
        p_wishbone_tx_fifo_fifo_7_18, p_wishbone_tx_fifo_fifo_7_19, 
        p_wishbone_tx_fifo_fifo_7_20, p_wishbone_tx_fifo_fifo_7_21, 
        p_wishbone_tx_fifo_fifo_7_22, p_wishbone_tx_fifo_fifo_7_23, 
        p_wishbone_tx_fifo_fifo_7_24, p_wishbone_tx_fifo_fifo_7_25, 
        p_wishbone_tx_fifo_fifo_7_26, p_wishbone_tx_fifo_fifo_7_27, 
        p_wishbone_tx_fifo_fifo_7_28, p_wishbone_tx_fifo_fifo_7_29, 
        p_wishbone_tx_fifo_fifo_7_30, p_wishbone_tx_fifo_fifo_7_31, 
        p_wishbone_tx_fifo_fifo_6_0, p_wishbone_tx_fifo_fifo_6_1, 
        p_wishbone_tx_fifo_fifo_6_2, p_wishbone_tx_fifo_fifo_6_3, 
        p_wishbone_tx_fifo_fifo_6_4, p_wishbone_tx_fifo_fifo_6_5, 
        p_wishbone_tx_fifo_fifo_6_6, p_wishbone_tx_fifo_fifo_6_7, 
        p_wishbone_tx_fifo_fifo_6_8, p_wishbone_tx_fifo_fifo_6_9, 
        p_wishbone_tx_fifo_fifo_6_10, p_wishbone_tx_fifo_fifo_6_11, 
        p_wishbone_tx_fifo_fifo_6_12, p_wishbone_tx_fifo_fifo_6_13, 
        p_wishbone_tx_fifo_fifo_6_14, p_wishbone_tx_fifo_fifo_6_15, 
        p_wishbone_tx_fifo_fifo_6_16, p_wishbone_tx_fifo_fifo_6_17, 
        p_wishbone_tx_fifo_fifo_6_18, p_wishbone_tx_fifo_fifo_6_19, 
        p_wishbone_tx_fifo_fifo_6_20, p_wishbone_tx_fifo_fifo_6_21, 
        p_wishbone_tx_fifo_fifo_6_22, p_wishbone_tx_fifo_fifo_6_23, 
        p_wishbone_tx_fifo_fifo_6_24, p_wishbone_tx_fifo_fifo_6_25, 
        p_wishbone_tx_fifo_fifo_6_26, p_wishbone_tx_fifo_fifo_6_27, 
        p_wishbone_tx_fifo_fifo_6_28, p_wishbone_tx_fifo_fifo_6_29, 
        p_wishbone_tx_fifo_fifo_6_30, p_wishbone_tx_fifo_fifo_6_31, 
        p_wishbone_tx_fifo_fifo_5_0, p_wishbone_tx_fifo_fifo_5_1, 
        p_wishbone_tx_fifo_fifo_5_2, p_wishbone_tx_fifo_fifo_5_3, 
        p_wishbone_tx_fifo_fifo_5_4, p_wishbone_tx_fifo_fifo_5_5, 
        p_wishbone_tx_fifo_fifo_5_6, p_wishbone_tx_fifo_fifo_5_7, 
        p_wishbone_tx_fifo_fifo_5_8, p_wishbone_tx_fifo_fifo_5_9, 
        p_wishbone_tx_fifo_fifo_5_10, p_wishbone_tx_fifo_fifo_5_11, 
        p_wishbone_tx_fifo_fifo_5_12, p_wishbone_tx_fifo_fifo_5_13, 
        p_wishbone_tx_fifo_fifo_5_14, p_wishbone_tx_fifo_fifo_5_15, 
        p_wishbone_tx_fifo_fifo_5_16, p_wishbone_tx_fifo_fifo_5_17, 
        p_wishbone_tx_fifo_fifo_5_18, p_wishbone_tx_fifo_fifo_5_19, 
        p_wishbone_tx_fifo_fifo_5_20, p_wishbone_tx_fifo_fifo_5_21, 
        p_wishbone_tx_fifo_fifo_5_22, p_wishbone_tx_fifo_fifo_5_23, 
        p_wishbone_tx_fifo_fifo_5_24, p_wishbone_tx_fifo_fifo_5_25, 
        p_wishbone_tx_fifo_fifo_5_26, p_wishbone_tx_fifo_fifo_5_27, 
        p_wishbone_tx_fifo_fifo_5_28, p_wishbone_tx_fifo_fifo_5_29, 
        p_wishbone_tx_fifo_fifo_5_30, p_wishbone_tx_fifo_fifo_5_31, 
        p_wishbone_tx_fifo_fifo_4_0, p_wishbone_tx_fifo_fifo_4_1, 
        p_wishbone_tx_fifo_fifo_4_2, p_wishbone_tx_fifo_fifo_4_3, 
        p_wishbone_tx_fifo_fifo_4_4, p_wishbone_tx_fifo_fifo_4_5, 
        p_wishbone_tx_fifo_fifo_4_6, p_wishbone_tx_fifo_fifo_4_7, 
        p_wishbone_tx_fifo_fifo_4_8, p_wishbone_tx_fifo_fifo_4_9, 
        p_wishbone_tx_fifo_fifo_4_10, p_wishbone_tx_fifo_fifo_4_11, 
        p_wishbone_tx_fifo_fifo_4_12, p_wishbone_tx_fifo_fifo_4_13, 
        p_wishbone_tx_fifo_fifo_4_14, p_wishbone_tx_fifo_fifo_4_15, 
        p_wishbone_tx_fifo_fifo_4_16, p_wishbone_tx_fifo_fifo_4_17, 
        p_wishbone_tx_fifo_fifo_4_18, p_wishbone_tx_fifo_fifo_4_19, 
        p_wishbone_tx_fifo_fifo_4_20, p_wishbone_tx_fifo_fifo_4_21, 
        p_wishbone_tx_fifo_fifo_4_22, p_wishbone_tx_fifo_fifo_4_23, 
        p_wishbone_tx_fifo_fifo_4_24, p_wishbone_tx_fifo_fifo_4_25, 
        p_wishbone_tx_fifo_fifo_4_26, p_wishbone_tx_fifo_fifo_4_27, 
        p_wishbone_tx_fifo_fifo_4_28, p_wishbone_tx_fifo_fifo_4_29, 
        p_wishbone_tx_fifo_fifo_4_30, p_wishbone_tx_fifo_fifo_4_31, 
        p_wishbone_tx_fifo_fifo_3_0, p_wishbone_tx_fifo_fifo_3_1, 
        p_wishbone_tx_fifo_fifo_3_2, p_wishbone_tx_fifo_fifo_3_3, 
        p_wishbone_tx_fifo_fifo_3_4, p_wishbone_tx_fifo_fifo_3_5, 
        p_wishbone_tx_fifo_fifo_3_6, p_wishbone_tx_fifo_fifo_3_7, 
        p_wishbone_tx_fifo_fifo_3_8, p_wishbone_tx_fifo_fifo_3_9, 
        p_wishbone_tx_fifo_fifo_3_10, p_wishbone_tx_fifo_fifo_3_11, 
        p_wishbone_tx_fifo_fifo_3_12, p_wishbone_tx_fifo_fifo_3_13, 
        p_wishbone_tx_fifo_fifo_3_14, p_wishbone_tx_fifo_fifo_3_15, 
        p_wishbone_tx_fifo_fifo_3_16, p_wishbone_tx_fifo_fifo_3_17, 
        p_wishbone_tx_fifo_fifo_3_18, p_wishbone_tx_fifo_fifo_3_19, 
        p_wishbone_tx_fifo_fifo_3_20, p_wishbone_tx_fifo_fifo_3_21, 
        p_wishbone_tx_fifo_fifo_3_22, p_wishbone_tx_fifo_fifo_3_23, 
        p_wishbone_tx_fifo_fifo_3_24, p_wishbone_tx_fifo_fifo_3_25, 
        p_wishbone_tx_fifo_fifo_3_26, p_wishbone_tx_fifo_fifo_3_27, 
        p_wishbone_tx_fifo_fifo_3_28, p_wishbone_tx_fifo_fifo_3_29, 
        p_wishbone_tx_fifo_fifo_3_30, p_wishbone_tx_fifo_fifo_3_31, 
        p_wishbone_tx_fifo_fifo_2_0, p_wishbone_tx_fifo_fifo_2_1, 
        p_wishbone_tx_fifo_fifo_2_2, p_wishbone_tx_fifo_fifo_2_3, 
        p_wishbone_tx_fifo_fifo_2_4, p_wishbone_tx_fifo_fifo_2_5, 
        p_wishbone_tx_fifo_fifo_2_6, p_wishbone_tx_fifo_fifo_2_7, 
        p_wishbone_tx_fifo_fifo_2_8, p_wishbone_tx_fifo_fifo_2_9, 
        p_wishbone_tx_fifo_fifo_2_10, p_wishbone_tx_fifo_fifo_2_11, 
        p_wishbone_tx_fifo_fifo_2_12, p_wishbone_tx_fifo_fifo_2_13, 
        p_wishbone_tx_fifo_fifo_2_14, p_wishbone_tx_fifo_fifo_2_15, 
        p_wishbone_tx_fifo_fifo_2_16, p_wishbone_tx_fifo_fifo_2_17, 
        p_wishbone_tx_fifo_fifo_2_18, p_wishbone_tx_fifo_fifo_2_19, 
        p_wishbone_tx_fifo_fifo_2_20, p_wishbone_tx_fifo_fifo_2_21, 
        p_wishbone_tx_fifo_fifo_2_22, p_wishbone_tx_fifo_fifo_2_23, 
        p_wishbone_tx_fifo_fifo_2_24, p_wishbone_tx_fifo_fifo_2_25, 
        p_wishbone_tx_fifo_fifo_2_26, p_wishbone_tx_fifo_fifo_2_27, 
        p_wishbone_tx_fifo_fifo_2_28, p_wishbone_tx_fifo_fifo_2_29, 
        p_wishbone_tx_fifo_fifo_2_30, p_wishbone_tx_fifo_fifo_2_31, 
        p_wishbone_tx_fifo_fifo_1_0, p_wishbone_tx_fifo_fifo_1_1, 
        p_wishbone_tx_fifo_fifo_1_2, p_wishbone_tx_fifo_fifo_1_3, 
        p_wishbone_tx_fifo_fifo_1_4, p_wishbone_tx_fifo_fifo_1_5, 
        p_wishbone_tx_fifo_fifo_1_6, p_wishbone_tx_fifo_fifo_1_7, 
        p_wishbone_tx_fifo_fifo_1_8, p_wishbone_tx_fifo_fifo_1_9, 
        p_wishbone_tx_fifo_fifo_1_10, p_wishbone_tx_fifo_fifo_1_11, 
        p_wishbone_tx_fifo_fifo_1_12, p_wishbone_tx_fifo_fifo_1_13, 
        p_wishbone_tx_fifo_fifo_1_14, p_wishbone_tx_fifo_fifo_1_15, 
        p_wishbone_tx_fifo_fifo_1_16, p_wishbone_tx_fifo_fifo_1_17, 
        p_wishbone_tx_fifo_fifo_1_18, p_wishbone_tx_fifo_fifo_1_19, 
        p_wishbone_tx_fifo_fifo_1_20, p_wishbone_tx_fifo_fifo_1_21, 
        p_wishbone_tx_fifo_fifo_1_22, p_wishbone_tx_fifo_fifo_1_23, 
        p_wishbone_tx_fifo_fifo_1_24, p_wishbone_tx_fifo_fifo_1_25, 
        p_wishbone_tx_fifo_fifo_1_26, p_wishbone_tx_fifo_fifo_1_27, 
        p_wishbone_tx_fifo_fifo_1_28, p_wishbone_tx_fifo_fifo_1_29, 
        p_wishbone_tx_fifo_fifo_1_30, p_wishbone_tx_fifo_fifo_1_31, 
        p_wishbone_tx_fifo_fifo_0_0, p_wishbone_tx_fifo_fifo_0_1, 
        p_wishbone_tx_fifo_fifo_0_2, p_wishbone_tx_fifo_fifo_0_3, 
        p_wishbone_tx_fifo_fifo_0_4, p_wishbone_tx_fifo_fifo_0_5, 
        p_wishbone_tx_fifo_fifo_0_6, p_wishbone_tx_fifo_fifo_0_7, 
        p_wishbone_tx_fifo_fifo_0_8, p_wishbone_tx_fifo_fifo_0_9, 
        p_wishbone_tx_fifo_fifo_0_10, p_wishbone_tx_fifo_fifo_0_11, 
        p_wishbone_tx_fifo_fifo_0_12, p_wishbone_tx_fifo_fifo_0_13, 
        p_wishbone_tx_fifo_fifo_0_14, p_wishbone_tx_fifo_fifo_0_15, 
        p_wishbone_tx_fifo_fifo_0_16, p_wishbone_tx_fifo_fifo_0_17, 
        p_wishbone_tx_fifo_fifo_0_18, p_wishbone_tx_fifo_fifo_0_19, 
        p_wishbone_tx_fifo_fifo_0_20, p_wishbone_tx_fifo_fifo_0_21, 
        p_wishbone_tx_fifo_fifo_0_22, p_wishbone_tx_fifo_fifo_0_23, 
        p_wishbone_tx_fifo_fifo_0_24, p_wishbone_tx_fifo_fifo_0_25, 
        p_wishbone_tx_fifo_fifo_0_26, p_wishbone_tx_fifo_fifo_0_27, 
        p_wishbone_tx_fifo_fifo_0_28, p_wishbone_tx_fifo_fifo_0_29, 
        p_wishbone_tx_fifo_fifo_0_30, p_wishbone_tx_fifo_fifo_0_31, 
        p_wishbone_tx_fifo_write_pointer_3, p_wishbone_tx_fifo_write_pointer_2, 
        p_wishbone_tx_fifo_write_pointer_1, p_wishbone_tx_fifo_write_pointer_0, 
        p_wishbone_tx_fifo_N17, p_wishbone_tx_fifo_N16, p_wishbone_tx_fifo_N15, 
        p_wishbone_tx_fifo_N14, p_wishbone_txfifo_cnt_4, 
        p_wishbone_txfifo_cnt_3, p_wishbone_txfifo_cnt_2, 
        p_wishbone_txfifo_cnt_1, p_wishbone_txfifo_cnt_0, r_TxPauseTV_8, 
        r_TxPauseTV_9, r_TxPauseTV_10, r_TxPauseTV_11, r_TxPauseTV_12, 
        r_TxPauseTV_13, r_TxPauseTV_14, r_TxPauseTV_15, r_TxPauseTV_0, 
        r_TxPauseTV_1, r_TxPauseTV_2, r_TxPauseTV_3, r_TxPauseTV_4, 
        r_TxPauseTV_5, r_TxPauseTV_6, r_TxPauseTV_7, r_HASH1_24, r_HASH1_25, 
        r_HASH1_26, r_HASH1_27, r_HASH1_28, r_HASH1_29, r_HASH1_30, r_HASH1_31, 
        r_HASH1_16, r_HASH1_17, r_HASH1_18, r_HASH1_19, r_HASH1_20, r_HASH1_21, 
        r_HASH1_22, r_HASH1_23, r_HASH1_8, r_HASH1_9, r_HASH1_10, r_HASH1_11, 
        r_HASH1_12, r_HASH1_13, r_HASH1_14, r_HASH1_15, r_HASH1_0, r_HASH1_1, 
        r_HASH1_2, r_HASH1_3, r_HASH1_4, r_HASH1_5, r_HASH1_6, r_HASH1_7, 
        r_HASH0_24, r_HASH0_25, r_HASH0_26, r_HASH0_27, r_HASH0_28, r_HASH0_29, 
        r_HASH0_30, r_HASH0_31, r_HASH0_16, r_HASH0_17, r_HASH0_18, r_HASH0_19, 
        r_HASH0_20, r_HASH0_21, r_HASH0_22, r_HASH0_23, r_HASH0_8, r_HASH0_9, 
        r_HASH0_10, r_HASH0_11, r_HASH0_12, r_HASH0_13, r_HASH0_14, r_HASH0_15, 
        r_HASH0_0, r_HASH0_1, r_HASH0_2, r_HASH0_3, r_HASH0_4, r_HASH0_5, 
        r_HASH0_6, r_HASH0_7, r_MAC_40, r_MAC_41, r_MAC_42, r_MAC_43, r_MAC_44, 
        r_MAC_45, r_MAC_46, r_MAC_47, r_MAC_32, r_MAC_33, r_MAC_34, r_MAC_35, 
        r_MAC_36, r_MAC_37, r_MAC_38, r_MAC_39, r_MAC_24, r_MAC_25, r_MAC_26, 
        r_MAC_27, r_MAC_28, r_MAC_29, r_MAC_30, r_MAC_31, r_MAC_16, r_MAC_17, 
        r_MAC_18, r_MAC_19, r_MAC_20, r_MAC_21, r_MAC_22, r_MAC_23, r_MAC_8, 
        r_MAC_9, r_MAC_10, r_MAC_11, r_MAC_12, r_MAC_13, r_MAC_14, r_MAC_15, 
        r_MAC_0, r_MAC_1, r_MAC_2, r_MAC_3, r_MAC_4, r_MAC_5, r_MAC_6, r_MAC_7, 
        r_CtrlData_8, r_CtrlData_9, r_CtrlData_10, r_CtrlData_11, 
        r_CtrlData_12, r_CtrlData_13, r_CtrlData_14, r_CtrlData_15, 
        r_CtrlData_0, r_CtrlData_1, r_CtrlData_2, r_CtrlData_3, r_CtrlData_4, 
        r_CtrlData_5, r_CtrlData_6, r_CtrlData_7, r_MinFL_8, r_MinFL_9, 
        r_MinFL_10, r_MinFL_11, r_MinFL_12, r_MinFL_13, r_MinFL_14, r_MinFL_15, 
        r_MaxFL_0, r_MaxFL_1, r_MaxFL_2, r_MaxFL_3, r_MaxFL_4, r_MaxFL_5, 
        r_MaxFL_6, r_MaxFL_7, r_TxPauseRq, r_MiiNoPre, r_IPGR2_0, r_IPGR2_1, 
        r_IPGR2_2, r_IPGR2_3, r_IPGR2_4, r_IPGR2_5, r_IPGR2_6, r_TxBDNum_0, 
        r_TxBDNum_1, r_TxBDNum_2, r_TxBDNum_3, r_TxBDNum_4, r_TxBDNum_5, 
        r_TxBDNum_6, r_TxBDNum_7, r_RGAD_0, r_RGAD_1, r_RGAD_2, r_RGAD_3, 
        r_RGAD_4, p_rxethmac1_crcrx_Crc_22, p_rxethmac1_crcrx_Crc_18, 
        p_rxethmac1_crcrx_Crc_14, p_rxethmac1_crcrx_Crc_10, 
        p_rxethmac1_crcrx_Crc_6, p_rxethmac1_crcrx_Crc_2, 
        p_rxethmac1_crcrx_Crc_5, p_rxethmac1_crcrx_Crc_23, 
        p_rxethmac1_crcrx_Crc_19, p_rxethmac1_crcrx_Crc_15, 
        p_rxethmac1_crcrx_Crc_11, p_rxethmac1_crcrx_Crc_7, 
        p_rxethmac1_crcrx_Crc_3, p_rxethmac1_Crc_31, p_rxethmac1_Crc_27, 
        p_rxethmac1_crcrx_Crc_1, p_rxethmac1_Crc_29, p_rxethmac1_crcrx_Crc_25, 
        p_rxethmac1_crcrx_Crc_21, p_rxethmac1_crcrx_Crc_17, 
        p_rxethmac1_crcrx_Crc_13, p_rxethmac1_crcrx_Crc_9, p_rxethmac1_Crc_30, 
        p_rxethmac1_Crc_26, p_rxethmac1_Crc_28, p_rxethmac1_crcrx_Crc_24, 
        p_rxethmac1_crcrx_Crc_20, p_rxethmac1_crcrx_Crc_16, 
        p_rxethmac1_crcrx_Crc_12, p_rxethmac1_crcrx_Crc_8, 
        p_rxethmac1_crcrx_Crc_4, p_rxethmac1_crcrx_Crc_0, 
        p_wishbone_rx_fifo_fifo_15_0, p_wishbone_rx_fifo_fifo_15_1, 
        p_wishbone_rx_fifo_fifo_15_2, p_wishbone_rx_fifo_fifo_15_3, 
        p_wishbone_rx_fifo_fifo_15_4, p_wishbone_rx_fifo_fifo_15_5, 
        p_wishbone_rx_fifo_fifo_15_6, p_wishbone_rx_fifo_fifo_15_7, 
        p_wishbone_rx_fifo_fifo_15_8, p_wishbone_rx_fifo_fifo_15_9, 
        p_wishbone_rx_fifo_fifo_15_10, p_wishbone_rx_fifo_fifo_15_11, 
        p_wishbone_rx_fifo_fifo_15_12, p_wishbone_rx_fifo_fifo_15_13, 
        p_wishbone_rx_fifo_fifo_15_14, p_wishbone_rx_fifo_fifo_15_15, 
        p_wishbone_rx_fifo_fifo_15_16, p_wishbone_rx_fifo_fifo_15_17, 
        p_wishbone_rx_fifo_fifo_15_18, p_wishbone_rx_fifo_fifo_15_19, 
        p_wishbone_rx_fifo_fifo_15_20, p_wishbone_rx_fifo_fifo_15_21, 
        p_wishbone_rx_fifo_fifo_15_22, p_wishbone_rx_fifo_fifo_15_23, 
        p_wishbone_rx_fifo_fifo_15_24, p_wishbone_rx_fifo_fifo_15_25, 
        p_wishbone_rx_fifo_fifo_15_26, p_wishbone_rx_fifo_fifo_15_27, 
        p_wishbone_rx_fifo_fifo_15_28, p_wishbone_rx_fifo_fifo_15_29, 
        p_wishbone_rx_fifo_fifo_15_30, p_wishbone_rx_fifo_fifo_15_31, 
        p_wishbone_rx_fifo_fifo_14_0, p_wishbone_rx_fifo_fifo_14_1, 
        p_wishbone_rx_fifo_fifo_14_2, p_wishbone_rx_fifo_fifo_14_3, 
        p_wishbone_rx_fifo_fifo_14_4, p_wishbone_rx_fifo_fifo_14_5, 
        p_wishbone_rx_fifo_fifo_14_6, p_wishbone_rx_fifo_fifo_14_7, 
        p_wishbone_rx_fifo_fifo_14_8, p_wishbone_rx_fifo_fifo_14_9, 
        p_wishbone_rx_fifo_fifo_14_10, p_wishbone_rx_fifo_fifo_14_11, 
        p_wishbone_rx_fifo_fifo_14_12, p_wishbone_rx_fifo_fifo_14_13, 
        p_wishbone_rx_fifo_fifo_14_14, p_wishbone_rx_fifo_fifo_14_15, 
        p_wishbone_rx_fifo_fifo_14_16, p_wishbone_rx_fifo_fifo_14_17, 
        p_wishbone_rx_fifo_fifo_14_18, p_wishbone_rx_fifo_fifo_14_19, 
        p_wishbone_rx_fifo_fifo_14_20, p_wishbone_rx_fifo_fifo_14_21, 
        p_wishbone_rx_fifo_fifo_14_22, p_wishbone_rx_fifo_fifo_14_23, 
        p_wishbone_rx_fifo_fifo_14_24, p_wishbone_rx_fifo_fifo_14_25, 
        p_wishbone_rx_fifo_fifo_14_26, p_wishbone_rx_fifo_fifo_14_27, 
        p_wishbone_rx_fifo_fifo_14_28, p_wishbone_rx_fifo_fifo_14_29, 
        p_wishbone_rx_fifo_fifo_14_30, p_wishbone_rx_fifo_fifo_14_31, 
        p_wishbone_rx_fifo_fifo_13_0, p_wishbone_rx_fifo_fifo_13_1, 
        p_wishbone_rx_fifo_fifo_13_2, p_wishbone_rx_fifo_fifo_13_3, 
        p_wishbone_rx_fifo_fifo_13_4, p_wishbone_rx_fifo_fifo_13_5, 
        p_wishbone_rx_fifo_fifo_13_6, p_wishbone_rx_fifo_fifo_13_7, 
        p_wishbone_rx_fifo_fifo_13_8, p_wishbone_rx_fifo_fifo_13_9, 
        p_wishbone_rx_fifo_fifo_13_10, p_wishbone_rx_fifo_fifo_13_11, 
        p_wishbone_rx_fifo_fifo_13_12, p_wishbone_rx_fifo_fifo_13_13, 
        p_wishbone_rx_fifo_fifo_13_14, p_wishbone_rx_fifo_fifo_13_15, 
        p_wishbone_rx_fifo_fifo_13_16, p_wishbone_rx_fifo_fifo_13_17, 
        p_wishbone_rx_fifo_fifo_13_18, p_wishbone_rx_fifo_fifo_13_19, 
        p_wishbone_rx_fifo_fifo_13_20, p_wishbone_rx_fifo_fifo_13_21, 
        p_wishbone_rx_fifo_fifo_13_22, p_wishbone_rx_fifo_fifo_13_23, 
        p_wishbone_rx_fifo_fifo_13_24, p_wishbone_rx_fifo_fifo_13_25, 
        p_wishbone_rx_fifo_fifo_13_26, p_wishbone_rx_fifo_fifo_13_27, 
        p_wishbone_rx_fifo_fifo_13_28, p_wishbone_rx_fifo_fifo_13_29, 
        p_wishbone_rx_fifo_fifo_13_30, p_wishbone_rx_fifo_fifo_13_31, 
        p_wishbone_rx_fifo_fifo_12_0, p_wishbone_rx_fifo_fifo_12_1, 
        p_wishbone_rx_fifo_fifo_12_2, p_wishbone_rx_fifo_fifo_12_3, 
        p_wishbone_rx_fifo_fifo_12_4, p_wishbone_rx_fifo_fifo_12_5, 
        p_wishbone_rx_fifo_fifo_12_6, p_wishbone_rx_fifo_fifo_12_7, 
        p_wishbone_rx_fifo_fifo_12_8, p_wishbone_rx_fifo_fifo_12_9, 
        p_wishbone_rx_fifo_fifo_12_10, p_wishbone_rx_fifo_fifo_12_11, 
        p_wishbone_rx_fifo_fifo_12_12, p_wishbone_rx_fifo_fifo_12_13, 
        p_wishbone_rx_fifo_fifo_12_14, p_wishbone_rx_fifo_fifo_12_15, 
        p_wishbone_rx_fifo_fifo_12_16, p_wishbone_rx_fifo_fifo_12_17, 
        p_wishbone_rx_fifo_fifo_12_18, p_wishbone_rx_fifo_fifo_12_19, 
        p_wishbone_rx_fifo_fifo_12_20, p_wishbone_rx_fifo_fifo_12_21, 
        p_wishbone_rx_fifo_fifo_12_22, p_wishbone_rx_fifo_fifo_12_23, 
        p_wishbone_rx_fifo_fifo_12_24, p_wishbone_rx_fifo_fifo_12_25, 
        p_wishbone_rx_fifo_fifo_12_26, p_wishbone_rx_fifo_fifo_12_27, 
        p_wishbone_rx_fifo_fifo_12_28, p_wishbone_rx_fifo_fifo_12_29, 
        p_wishbone_rx_fifo_fifo_12_30, p_wishbone_rx_fifo_fifo_12_31, 
        p_wishbone_rx_fifo_fifo_11_0, p_wishbone_rx_fifo_fifo_11_1, 
        p_wishbone_rx_fifo_fifo_11_2, p_wishbone_rx_fifo_fifo_11_3, 
        p_wishbone_rx_fifo_fifo_11_4, p_wishbone_rx_fifo_fifo_11_5, 
        p_wishbone_rx_fifo_fifo_11_6, p_wishbone_rx_fifo_fifo_11_7, 
        p_wishbone_rx_fifo_fifo_11_8, p_wishbone_rx_fifo_fifo_11_9, 
        p_wishbone_rx_fifo_fifo_11_10, p_wishbone_rx_fifo_fifo_11_11, 
        p_wishbone_rx_fifo_fifo_11_12, p_wishbone_rx_fifo_fifo_11_13, 
        p_wishbone_rx_fifo_fifo_11_14, p_wishbone_rx_fifo_fifo_11_15, 
        p_wishbone_rx_fifo_fifo_11_16, p_wishbone_rx_fifo_fifo_11_17, 
        p_wishbone_rx_fifo_fifo_11_18, p_wishbone_rx_fifo_fifo_11_19, 
        p_wishbone_rx_fifo_fifo_11_20, p_wishbone_rx_fifo_fifo_11_21, 
        p_wishbone_rx_fifo_fifo_11_22, p_wishbone_rx_fifo_fifo_11_23, 
        p_wishbone_rx_fifo_fifo_11_24, p_wishbone_rx_fifo_fifo_11_25, 
        p_wishbone_rx_fifo_fifo_11_26, p_wishbone_rx_fifo_fifo_11_27, 
        p_wishbone_rx_fifo_fifo_11_28, p_wishbone_rx_fifo_fifo_11_29, 
        p_wishbone_rx_fifo_fifo_11_30, p_wishbone_rx_fifo_fifo_11_31, 
        p_wishbone_rx_fifo_fifo_10_0, p_wishbone_rx_fifo_fifo_10_1, 
        p_wishbone_rx_fifo_fifo_10_2, p_wishbone_rx_fifo_fifo_10_3, 
        p_wishbone_rx_fifo_fifo_10_4, p_wishbone_rx_fifo_fifo_10_5, 
        p_wishbone_rx_fifo_fifo_10_6, p_wishbone_rx_fifo_fifo_10_7, 
        p_wishbone_rx_fifo_fifo_10_8, p_wishbone_rx_fifo_fifo_10_9, 
        p_wishbone_rx_fifo_fifo_10_10, p_wishbone_rx_fifo_fifo_10_11, 
        p_wishbone_rx_fifo_fifo_10_12, p_wishbone_rx_fifo_fifo_10_13, 
        p_wishbone_rx_fifo_fifo_10_14, p_wishbone_rx_fifo_fifo_10_15, 
        p_wishbone_rx_fifo_fifo_10_16, p_wishbone_rx_fifo_fifo_10_17, 
        p_wishbone_rx_fifo_fifo_10_18, p_wishbone_rx_fifo_fifo_10_19, 
        p_wishbone_rx_fifo_fifo_10_20, p_wishbone_rx_fifo_fifo_10_21, 
        p_wishbone_rx_fifo_fifo_10_22, p_wishbone_rx_fifo_fifo_10_23, 
        p_wishbone_rx_fifo_fifo_10_24, p_wishbone_rx_fifo_fifo_10_25, 
        p_wishbone_rx_fifo_fifo_10_26, p_wishbone_rx_fifo_fifo_10_27, 
        p_wishbone_rx_fifo_fifo_10_28, p_wishbone_rx_fifo_fifo_10_29, 
        p_wishbone_rx_fifo_fifo_10_30, p_wishbone_rx_fifo_fifo_10_31, 
        p_wishbone_rx_fifo_fifo_9_0, p_wishbone_rx_fifo_fifo_9_1, 
        p_wishbone_rx_fifo_fifo_9_2, p_wishbone_rx_fifo_fifo_9_3, 
        p_wishbone_rx_fifo_fifo_9_4, p_wishbone_rx_fifo_fifo_9_5, 
        p_wishbone_rx_fifo_fifo_9_6, p_wishbone_rx_fifo_fifo_9_7, 
        p_wishbone_rx_fifo_fifo_9_8, p_wishbone_rx_fifo_fifo_9_9, 
        p_wishbone_rx_fifo_fifo_9_10, p_wishbone_rx_fifo_fifo_9_11, 
        p_wishbone_rx_fifo_fifo_9_12, p_wishbone_rx_fifo_fifo_9_13, 
        p_wishbone_rx_fifo_fifo_9_14, p_wishbone_rx_fifo_fifo_9_15, 
        p_wishbone_rx_fifo_fifo_9_16, p_wishbone_rx_fifo_fifo_9_17, 
        p_wishbone_rx_fifo_fifo_9_18, p_wishbone_rx_fifo_fifo_9_19, 
        p_wishbone_rx_fifo_fifo_9_20, p_wishbone_rx_fifo_fifo_9_21, 
        p_wishbone_rx_fifo_fifo_9_22, p_wishbone_rx_fifo_fifo_9_23, 
        p_wishbone_rx_fifo_fifo_9_24, p_wishbone_rx_fifo_fifo_9_25, 
        p_wishbone_rx_fifo_fifo_9_26, p_wishbone_rx_fifo_fifo_9_27, 
        p_wishbone_rx_fifo_fifo_9_28, p_wishbone_rx_fifo_fifo_9_29, 
        p_wishbone_rx_fifo_fifo_9_30, p_wishbone_rx_fifo_fifo_9_31, 
        p_wishbone_rx_fifo_fifo_8_0, p_wishbone_rx_fifo_fifo_8_1, 
        p_wishbone_rx_fifo_fifo_8_2, p_wishbone_rx_fifo_fifo_8_3, 
        p_wishbone_rx_fifo_fifo_8_4, p_wishbone_rx_fifo_fifo_8_5, 
        p_wishbone_rx_fifo_fifo_8_6, p_wishbone_rx_fifo_fifo_8_7, 
        p_wishbone_rx_fifo_fifo_8_8, p_wishbone_rx_fifo_fifo_8_9, 
        p_wishbone_rx_fifo_fifo_8_10, p_wishbone_rx_fifo_fifo_8_11, 
        p_wishbone_rx_fifo_fifo_8_12, p_wishbone_rx_fifo_fifo_8_13, 
        p_wishbone_rx_fifo_fifo_8_14, p_wishbone_rx_fifo_fifo_8_15, 
        p_wishbone_rx_fifo_fifo_8_16, p_wishbone_rx_fifo_fifo_8_17, 
        p_wishbone_rx_fifo_fifo_8_18, p_wishbone_rx_fifo_fifo_8_19, 
        p_wishbone_rx_fifo_fifo_8_20, p_wishbone_rx_fifo_fifo_8_21, 
        p_wishbone_rx_fifo_fifo_8_22, p_wishbone_rx_fifo_fifo_8_23, 
        p_wishbone_rx_fifo_fifo_8_24, p_wishbone_rx_fifo_fifo_8_25, 
        p_wishbone_rx_fifo_fifo_8_26, p_wishbone_rx_fifo_fifo_8_27, 
        p_wishbone_rx_fifo_fifo_8_28, p_wishbone_rx_fifo_fifo_8_29, 
        p_wishbone_rx_fifo_fifo_8_30, p_wishbone_rx_fifo_fifo_8_31, 
        p_wishbone_rx_fifo_fifo_7_0, p_wishbone_rx_fifo_fifo_7_1, 
        p_wishbone_rx_fifo_fifo_7_2, p_wishbone_rx_fifo_fifo_7_3, 
        p_wishbone_rx_fifo_fifo_7_4, p_wishbone_rx_fifo_fifo_7_5, 
        p_wishbone_rx_fifo_fifo_7_6, p_wishbone_rx_fifo_fifo_7_7, 
        p_wishbone_rx_fifo_fifo_7_8, p_wishbone_rx_fifo_fifo_7_9, 
        p_wishbone_rx_fifo_fifo_7_10, p_wishbone_rx_fifo_fifo_7_11, 
        p_wishbone_rx_fifo_fifo_7_12, p_wishbone_rx_fifo_fifo_7_13, 
        p_wishbone_rx_fifo_fifo_7_14, p_wishbone_rx_fifo_fifo_7_15, 
        p_wishbone_rx_fifo_fifo_7_16, p_wishbone_rx_fifo_fifo_7_17, 
        p_wishbone_rx_fifo_fifo_7_18, p_wishbone_rx_fifo_fifo_7_19, 
        p_wishbone_rx_fifo_fifo_7_20, p_wishbone_rx_fifo_fifo_7_21, 
        p_wishbone_rx_fifo_fifo_7_22, p_wishbone_rx_fifo_fifo_7_23, 
        p_wishbone_rx_fifo_fifo_7_24, p_wishbone_rx_fifo_fifo_7_25, 
        p_wishbone_rx_fifo_fifo_7_26, p_wishbone_rx_fifo_fifo_7_27, 
        p_wishbone_rx_fifo_fifo_7_28, p_wishbone_rx_fifo_fifo_7_29, 
        p_wishbone_rx_fifo_fifo_7_30, p_wishbone_rx_fifo_fifo_7_31, 
        p_wishbone_rx_fifo_fifo_6_0, p_wishbone_rx_fifo_fifo_6_1, 
        p_wishbone_rx_fifo_fifo_6_2, p_wishbone_rx_fifo_fifo_6_3, 
        p_wishbone_rx_fifo_fifo_6_4, p_wishbone_rx_fifo_fifo_6_5, 
        p_wishbone_rx_fifo_fifo_6_6, p_wishbone_rx_fifo_fifo_6_7, 
        p_wishbone_rx_fifo_fifo_6_8, p_wishbone_rx_fifo_fifo_6_9, 
        p_wishbone_rx_fifo_fifo_6_10, p_wishbone_rx_fifo_fifo_6_11, 
        p_wishbone_rx_fifo_fifo_6_12, p_wishbone_rx_fifo_fifo_6_13, 
        p_wishbone_rx_fifo_fifo_6_14, p_wishbone_rx_fifo_fifo_6_15, 
        p_wishbone_rx_fifo_fifo_6_16, p_wishbone_rx_fifo_fifo_6_17, 
        p_wishbone_rx_fifo_fifo_6_18, p_wishbone_rx_fifo_fifo_6_19, 
        p_wishbone_rx_fifo_fifo_6_20, p_wishbone_rx_fifo_fifo_6_21, 
        p_wishbone_rx_fifo_fifo_6_22, p_wishbone_rx_fifo_fifo_6_23, 
        p_wishbone_rx_fifo_fifo_6_24, p_wishbone_rx_fifo_fifo_6_25, 
        p_wishbone_rx_fifo_fifo_6_26, p_wishbone_rx_fifo_fifo_6_27, 
        p_wishbone_rx_fifo_fifo_6_28, p_wishbone_rx_fifo_fifo_6_29, 
        p_wishbone_rx_fifo_fifo_6_30, p_wishbone_rx_fifo_fifo_6_31, 
        p_wishbone_rx_fifo_fifo_5_0, p_wishbone_rx_fifo_fifo_5_1, 
        p_wishbone_rx_fifo_fifo_5_2, p_wishbone_rx_fifo_fifo_5_3, 
        p_wishbone_rx_fifo_fifo_5_4, p_wishbone_rx_fifo_fifo_5_5, 
        p_wishbone_rx_fifo_fifo_5_6, p_wishbone_rx_fifo_fifo_5_7, 
        p_wishbone_rx_fifo_fifo_5_8, p_wishbone_rx_fifo_fifo_5_9, 
        p_wishbone_rx_fifo_fifo_5_10, p_wishbone_rx_fifo_fifo_5_11, 
        p_wishbone_rx_fifo_fifo_5_12, p_wishbone_rx_fifo_fifo_5_13, 
        p_wishbone_rx_fifo_fifo_5_14, p_wishbone_rx_fifo_fifo_5_15, 
        p_wishbone_rx_fifo_fifo_5_16, p_wishbone_rx_fifo_fifo_5_17, 
        p_wishbone_rx_fifo_fifo_5_18, p_wishbone_rx_fifo_fifo_5_19, 
        p_wishbone_rx_fifo_fifo_5_20, p_wishbone_rx_fifo_fifo_5_21, 
        p_wishbone_rx_fifo_fifo_5_22, p_wishbone_rx_fifo_fifo_5_23, 
        p_wishbone_rx_fifo_fifo_5_24, p_wishbone_rx_fifo_fifo_5_25, 
        p_wishbone_rx_fifo_fifo_5_26, p_wishbone_rx_fifo_fifo_5_27, 
        p_wishbone_rx_fifo_fifo_5_28, p_wishbone_rx_fifo_fifo_5_29, 
        p_wishbone_rx_fifo_fifo_5_30, p_wishbone_rx_fifo_fifo_5_31, 
        p_wishbone_rx_fifo_fifo_4_0, p_wishbone_rx_fifo_fifo_4_1, 
        p_wishbone_rx_fifo_fifo_4_2, p_wishbone_rx_fifo_fifo_4_3, 
        p_wishbone_rx_fifo_fifo_4_4, p_wishbone_rx_fifo_fifo_4_5, 
        p_wishbone_rx_fifo_fifo_4_6, p_wishbone_rx_fifo_fifo_4_7, 
        p_wishbone_rx_fifo_fifo_4_8, p_wishbone_rx_fifo_fifo_4_9, 
        p_wishbone_rx_fifo_fifo_4_10, p_wishbone_rx_fifo_fifo_4_11, 
        p_wishbone_rx_fifo_fifo_4_12, p_wishbone_rx_fifo_fifo_4_13, 
        p_wishbone_rx_fifo_fifo_4_14, p_wishbone_rx_fifo_fifo_4_15, 
        p_wishbone_rx_fifo_fifo_4_16, p_wishbone_rx_fifo_fifo_4_17, 
        p_wishbone_rx_fifo_fifo_4_18, p_wishbone_rx_fifo_fifo_4_19, 
        p_wishbone_rx_fifo_fifo_4_20, p_wishbone_rx_fifo_fifo_4_21, 
        p_wishbone_rx_fifo_fifo_4_22, p_wishbone_rx_fifo_fifo_4_23, 
        p_wishbone_rx_fifo_fifo_4_24, p_wishbone_rx_fifo_fifo_4_25, 
        p_wishbone_rx_fifo_fifo_4_26, p_wishbone_rx_fifo_fifo_4_27, 
        p_wishbone_rx_fifo_fifo_4_28, p_wishbone_rx_fifo_fifo_4_29, 
        p_wishbone_rx_fifo_fifo_4_30, p_wishbone_rx_fifo_fifo_4_31, 
        p_wishbone_rx_fifo_fifo_3_0, p_wishbone_rx_fifo_fifo_3_1, 
        p_wishbone_rx_fifo_fifo_3_2, p_wishbone_rx_fifo_fifo_3_3, 
        p_wishbone_rx_fifo_fifo_3_4, p_wishbone_rx_fifo_fifo_3_5, 
        p_wishbone_rx_fifo_fifo_3_6, p_wishbone_rx_fifo_fifo_3_7, 
        p_wishbone_rx_fifo_fifo_3_8, p_wishbone_rx_fifo_fifo_3_9, 
        p_wishbone_rx_fifo_fifo_3_10, p_wishbone_rx_fifo_fifo_3_11, 
        p_wishbone_rx_fifo_fifo_3_12, p_wishbone_rx_fifo_fifo_3_13, 
        p_wishbone_rx_fifo_fifo_3_14, p_wishbone_rx_fifo_fifo_3_15, 
        p_wishbone_rx_fifo_fifo_3_16, p_wishbone_rx_fifo_fifo_3_17, 
        p_wishbone_rx_fifo_fifo_3_18, p_wishbone_rx_fifo_fifo_3_19, 
        p_wishbone_rx_fifo_fifo_3_20, p_wishbone_rx_fifo_fifo_3_21, 
        p_wishbone_rx_fifo_fifo_3_22, p_wishbone_rx_fifo_fifo_3_23, 
        p_wishbone_rx_fifo_fifo_3_24, p_wishbone_rx_fifo_fifo_3_25, 
        p_wishbone_rx_fifo_fifo_3_26, p_wishbone_rx_fifo_fifo_3_27, 
        p_wishbone_rx_fifo_fifo_3_28, p_wishbone_rx_fifo_fifo_3_29, 
        p_wishbone_rx_fifo_fifo_3_30, p_wishbone_rx_fifo_fifo_3_31, 
        p_wishbone_rx_fifo_fifo_2_0, p_wishbone_rx_fifo_fifo_2_1, 
        p_wishbone_rx_fifo_fifo_2_2, p_wishbone_rx_fifo_fifo_2_3, 
        p_wishbone_rx_fifo_fifo_2_4, p_wishbone_rx_fifo_fifo_2_5, 
        p_wishbone_rx_fifo_fifo_2_6, p_wishbone_rx_fifo_fifo_2_7, 
        p_wishbone_rx_fifo_fifo_2_8, p_wishbone_rx_fifo_fifo_2_9, 
        p_wishbone_rx_fifo_fifo_2_10, p_wishbone_rx_fifo_fifo_2_11, 
        p_wishbone_rx_fifo_fifo_2_12, p_wishbone_rx_fifo_fifo_2_13, 
        p_wishbone_rx_fifo_fifo_2_14, p_wishbone_rx_fifo_fifo_2_15, 
        p_wishbone_rx_fifo_fifo_2_16, p_wishbone_rx_fifo_fifo_2_17, 
        p_wishbone_rx_fifo_fifo_2_18, p_wishbone_rx_fifo_fifo_2_19, 
        p_wishbone_rx_fifo_fifo_2_20, p_wishbone_rx_fifo_fifo_2_21, 
        p_wishbone_rx_fifo_fifo_2_22, p_wishbone_rx_fifo_fifo_2_23, 
        p_wishbone_rx_fifo_fifo_2_24, p_wishbone_rx_fifo_fifo_2_25, 
        p_wishbone_rx_fifo_fifo_2_26, p_wishbone_rx_fifo_fifo_2_27, 
        p_wishbone_rx_fifo_fifo_2_28, p_wishbone_rx_fifo_fifo_2_29, 
        p_wishbone_rx_fifo_fifo_2_30, p_wishbone_rx_fifo_fifo_2_31, 
        p_wishbone_rx_fifo_fifo_1_0, p_wishbone_rx_fifo_fifo_1_1, 
        p_wishbone_rx_fifo_fifo_1_2, p_wishbone_rx_fifo_fifo_1_3, 
        p_wishbone_rx_fifo_fifo_1_4, p_wishbone_rx_fifo_fifo_1_5, 
        p_wishbone_rx_fifo_fifo_1_6, p_wishbone_rx_fifo_fifo_1_7, 
        p_wishbone_rx_fifo_fifo_1_8, p_wishbone_rx_fifo_fifo_1_9, 
        p_wishbone_rx_fifo_fifo_1_10, p_wishbone_rx_fifo_fifo_1_11, 
        p_wishbone_rx_fifo_fifo_1_12, p_wishbone_rx_fifo_fifo_1_13, 
        p_wishbone_rx_fifo_fifo_1_14, p_wishbone_rx_fifo_fifo_1_15, 
        p_wishbone_rx_fifo_fifo_1_16, p_wishbone_rx_fifo_fifo_1_17, 
        p_wishbone_rx_fifo_fifo_1_18, p_wishbone_rx_fifo_fifo_1_19, 
        p_wishbone_rx_fifo_fifo_1_20, p_wishbone_rx_fifo_fifo_1_21, 
        p_wishbone_rx_fifo_fifo_1_22, p_wishbone_rx_fifo_fifo_1_23, 
        p_wishbone_rx_fifo_fifo_1_24, p_wishbone_rx_fifo_fifo_1_25, 
        p_wishbone_rx_fifo_fifo_1_26, p_wishbone_rx_fifo_fifo_1_27, 
        p_wishbone_rx_fifo_fifo_1_28, p_wishbone_rx_fifo_fifo_1_29, 
        p_wishbone_rx_fifo_fifo_1_30, p_wishbone_rx_fifo_fifo_1_31, 
        p_wishbone_rx_fifo_fifo_0_0, p_wishbone_rx_fifo_fifo_0_1, 
        p_wishbone_rx_fifo_fifo_0_2, p_wishbone_rx_fifo_fifo_0_3, 
        p_wishbone_rx_fifo_fifo_0_4, p_wishbone_rx_fifo_fifo_0_5, 
        p_wishbone_rx_fifo_fifo_0_6, p_wishbone_rx_fifo_fifo_0_7, 
        p_wishbone_rx_fifo_fifo_0_8, p_wishbone_rx_fifo_fifo_0_9, 
        p_wishbone_rx_fifo_fifo_0_10, p_wishbone_rx_fifo_fifo_0_11, 
        p_wishbone_rx_fifo_fifo_0_12, p_wishbone_rx_fifo_fifo_0_13, 
        p_wishbone_rx_fifo_fifo_0_14, p_wishbone_rx_fifo_fifo_0_15, 
        p_wishbone_rx_fifo_fifo_0_16, p_wishbone_rx_fifo_fifo_0_17, 
        p_wishbone_rx_fifo_fifo_0_18, p_wishbone_rx_fifo_fifo_0_19, 
        p_wishbone_rx_fifo_fifo_0_20, p_wishbone_rx_fifo_fifo_0_21, 
        p_wishbone_rx_fifo_fifo_0_22, p_wishbone_rx_fifo_fifo_0_23, 
        p_wishbone_rx_fifo_fifo_0_24, p_wishbone_rx_fifo_fifo_0_25, 
        p_wishbone_rx_fifo_fifo_0_26, p_wishbone_rx_fifo_fifo_0_27, 
        p_wishbone_rx_fifo_fifo_0_28, p_wishbone_rx_fifo_fifo_0_29, 
        p_wishbone_rx_fifo_fifo_0_30, p_wishbone_rx_fifo_fifo_0_31, 
        p_wishbone_rx_fifo_write_pointer_3, p_wishbone_rx_fifo_write_pointer_2, 
        p_wishbone_rx_fifo_write_pointer_1, p_wishbone_rx_fifo_write_pointer_0, 
        p_wishbone_rx_fifo_N17, p_wishbone_rx_fifo_N16, p_wishbone_rx_fifo_N15, 
        p_wishbone_rx_fifo_N14, p_wishbone_rxfifo_cnt_4, 
        p_wishbone_rxfifo_cnt_3, p_wishbone_rxfifo_cnt_2, 
        p_wishbone_rxfifo_cnt_1, p_wishbone_rxfifo_cnt_0, wb_dat_o_0, 
        wb_dat_o_1, wb_dat_o_2, wb_dat_o_3, wb_dat_o_4, wb_dat_o_5, wb_dat_o_6, 
        wb_dat_o_7, wb_dat_o_8, wb_dat_o_9, wb_dat_o_10, wb_dat_o_11, 
        wb_dat_o_12, wb_dat_o_13, wb_dat_o_14, wb_dat_o_15, wb_dat_o_16, 
        wb_dat_o_17, wb_dat_o_18, wb_dat_o_19, wb_dat_o_20, wb_dat_o_21, 
        wb_dat_o_22, wb_dat_o_23, wb_dat_o_24, wb_dat_o_25, wb_dat_o_26, 
        wb_dat_o_27, wb_dat_o_28, wb_dat_o_29, wb_dat_o_30, wb_dat_o_31, 
        m_wb_adr_o_0, m_wb_adr_o_1, m_wb_adr_o_2, m_wb_adr_o_3, m_wb_adr_o_4, 
        m_wb_adr_o_5, m_wb_adr_o_6, m_wb_adr_o_7, m_wb_adr_o_8, m_wb_adr_o_9, 
        m_wb_adr_o_10, m_wb_adr_o_11, m_wb_adr_o_12, m_wb_adr_o_13, 
        m_wb_adr_o_14, m_wb_adr_o_15, m_wb_adr_o_16, m_wb_adr_o_17, 
        m_wb_adr_o_18, m_wb_adr_o_19, m_wb_adr_o_20, m_wb_adr_o_21, 
        m_wb_adr_o_22, m_wb_adr_o_23, m_wb_adr_o_24, m_wb_adr_o_25, 
        m_wb_adr_o_26, m_wb_adr_o_27, m_wb_adr_o_28, m_wb_adr_o_29, 
        m_wb_adr_o_30, m_wb_adr_o_31, m_wb_sel_o_0, m_wb_sel_o_1, m_wb_sel_o_2, 
        m_wb_sel_o_3, m_wb_dat_o_0, m_wb_dat_o_1, m_wb_dat_o_2, m_wb_dat_o_3, 
        m_wb_dat_o_4, m_wb_dat_o_5, m_wb_dat_o_6, m_wb_dat_o_7, m_wb_dat_o_8, 
        m_wb_dat_o_9, m_wb_dat_o_10, m_wb_dat_o_11, m_wb_dat_o_12, 
        m_wb_dat_o_13, m_wb_dat_o_14, m_wb_dat_o_15, m_wb_dat_o_16, 
        m_wb_dat_o_17, m_wb_dat_o_18, m_wb_dat_o_19, m_wb_dat_o_20, 
        m_wb_dat_o_21, m_wb_dat_o_22, m_wb_dat_o_23, m_wb_dat_o_24, 
        m_wb_dat_o_25, m_wb_dat_o_26, m_wb_dat_o_27, m_wb_dat_o_28, 
        m_wb_dat_o_29, m_wb_dat_o_30, m_wb_dat_o_31, mtxd_pad_o_0, 
        mtxd_pad_o_1, mtxd_pad_o_2, mtxd_pad_o_3, wb_ack_o, wb_err_o, 
        m_wb_we_o, m_wb_cyc_o, m_wb_stb_o, mtxen_pad_o, mtxerr_pad_o, 
        mdc_pad_o, md_pad_o, md_padoe_o, int_o, N10, RxAbortRst_sync1, n126, 
        WillSendControlFrame, N23, N24, N25, n124, n125, WillTransmit, N9, 
        temp_wb_dat_o_0, temp_wb_dat_o_1, temp_wb_dat_o_2, temp_wb_dat_o_3, 
        temp_wb_dat_o_4, temp_wb_dat_o_5, temp_wb_dat_o_6, temp_wb_dat_o_7, 
        temp_wb_dat_o_8, temp_wb_dat_o_9, temp_wb_dat_o_10, temp_wb_dat_o_11, 
        temp_wb_dat_o_12, temp_wb_dat_o_13, temp_wb_dat_o_14, temp_wb_dat_o_15, 
        temp_wb_dat_o_16, temp_wb_dat_o_17, temp_wb_dat_o_18, temp_wb_dat_o_19, 
        temp_wb_dat_o_20, temp_wb_dat_o_21, temp_wb_dat_o_22, temp_wb_dat_o_23, 
        temp_wb_dat_o_24, temp_wb_dat_o_25, temp_wb_dat_o_26, temp_wb_dat_o_27, 
        temp_wb_dat_o_28, temp_wb_dat_o_29, temp_wb_dat_o_30, temp_wb_dat_o_31, 
        p_miim1_n133, p_miim1_n134, p_miim1_n135, p_miim1_n136, p_miim1_n153, 
        p_miim1_n137, p_miim1_n138, p_miim1_n139, p_miim1_n140, p_miim1_n141, 
        p_miim1_n142, p_miim1_n156, p_miim1_N9, p_miim1_n143, p_miim1_n144, 
        p_miim1_n145, p_miim1_n154, p_miim1_n146, p_miim1_n147, p_miim1_n155, 
        p_miim1_EndBusy_d, p_miim1_N8, p_miim1_n148, p_miim1_n149, 
        p_miim1_n150, p_miim1_n157, p_miim1_n151, p_miim1_WCtrlData_q2, 
        p_miim1_WCtrlData_q1, r_WCtrlData, p_miim1_RStat_q2, p_miim1_RStat_q1, 
        r_RStat, p_miim1_n152, p_miim1_ScanStat_q1, r_ScanStat, p_ethreg1_n678, 
        p_ethreg1_n679, p_ethreg1_n680, p_ethreg1_n681, p_ethreg1_n682, 
        p_ethreg1_n683, p_ethreg1_n684, p_ethreg1_N228, 
        p_ethreg1_ResetRxCIrq_sync1, p_ethreg1_SetRxCIrq_sync2, 
        p_ethreg1_SetRxCIrq_sync1, p_ethreg1_SetRxCIrq_rxclk, p_ethreg1_n685, 
        p_ethreg1_N222, p_ethreg1_SetTxCIrq_sync2, p_ethreg1_SetTxCIrq_sync1, 
        p_ethreg1_SetTxCIrq_txclk, p_ethreg1_n686, p_maccontrol1_n53, 
        p_maccontrol1_n54, TxDoneIn, TxAbortIn, p_maccontrol1_n55, 
        p_txethmac1_n152, p_txethmac1_n153, p_txethmac1_n149, 
        p_txethmac1_PacketFinished_d, p_txethmac1_n148, p_txethmac1_n147, 
        p_txethmac1_n150, p_txethmac1_n155, p_txethmac1_MTxD_d_0, 
        p_txethmac1_MTxD_d_1, p_txethmac1_MTxD_d_2, p_txethmac1_MTxD_d_3, 
        p_txethmac1_N88, p_txethmac1_N86, p_txethmac1_N87, p_txethmac1_n156, 
        p_txethmac1_N29, p_txethmac1_n151, p_txethmac1_n154, p_rxethmac1_n95, 
        p_rxethmac1_n94, p_rxethmac1_N51, p_rxethmac1_GenerateRxEndFrm, 
        p_rxethmac1_RxStartFrm_d, p_rxethmac1_GenerateRxStartFrm, 
        p_rxethmac1_RxValid_d, n33940, p_rxethmac1_RxData_d_7, 
        p_rxethmac1_n103, p_rxethmac1_RxData_d_6, p_rxethmac1_n102, 
        p_rxethmac1_RxData_d_5, p_rxethmac1_n101, p_rxethmac1_RxData_d_4, 
        p_rxethmac1_n100, p_rxethmac1_RxData_d_3, p_rxethmac1_n99, 
        p_rxethmac1_RxData_d_2, p_rxethmac1_n98, p_rxethmac1_RxData_d_1, 
        p_rxethmac1_n97, p_rxethmac1_RxData_d_0, p_rxethmac1_n96, 
        RxStateData_0, p_rxethmac1_LatchedByte_4, p_rxethmac1_LatchedByte_5, 
        p_rxethmac1_LatchedByte_6, p_rxethmac1_LatchedByte_7, MRxD_Lb_0, 
        MRxD_Lb_1, MRxD_Lb_2, MRxD_Lb_3, p_rxethmac1_n104, p_rxethmac1_n105, 
        p_rxethmac1_n106, p_rxethmac1_n107, p_rxethmac1_n108, p_rxethmac1_n109, 
        p_rxethmac1_N3, p_wishbone_Busy_IRQ_sync2, p_wishbone_Busy_IRQ_sync1, 
        p_wishbone_Busy_IRQ_rck, p_wishbone_n2138, p_wishbone_N1329, 
        p_wishbone_N1326, p_wishbone_N1322, p_wishbone_N1319, 
        RxStatusWriteLatched_sync2, p_wishbone_RxStatusWriteLatched_sync1, 
        p_wishbone_RxStatusWriteLatched, p_wishbone_n2139, p_wishbone_n2141, 
        p_wishbone_n2142, p_wishbone_n2143, p_wishbone_n2144, p_wishbone_n2145, 
        p_wishbone_n2146, p_wishbone_n2147, p_wishbone_n2148, p_wishbone_n2149, 
        p_wishbone_n2150, p_wishbone_n2151, p_wishbone_n2152, p_wishbone_n2153, 
        p_wishbone_n2154, p_wishbone_n2155, p_wishbone_n2156, p_wishbone_n2157, 
        p_wishbone_n2158, p_wishbone_n2159, p_wishbone_n2160, p_wishbone_n2161, 
        p_wishbone_n2162, p_wishbone_n2163, p_wishbone_n2164, p_wishbone_n2165, 
        p_wishbone_n2166, p_wishbone_n2167, p_wishbone_n2168, p_wishbone_n2169, 
        p_wishbone_n2140, p_wishbone_n2171, p_wishbone_n2172, p_wishbone_n2173, 
        p_wishbone_n2174, p_wishbone_n2175, p_wishbone_n2176, p_wishbone_n2177, 
        p_wishbone_n2178, p_wishbone_n2179, p_wishbone_n2180, p_wishbone_n2181, 
        p_wishbone_n2182, p_wishbone_n2183, p_wishbone_n2184, p_wishbone_n2185, 
        p_wishbone_n2186, p_wishbone_n2187, p_wishbone_n2188, p_wishbone_n2189, 
        p_wishbone_n2190, p_wishbone_n2191, p_wishbone_n2192, p_wishbone_n2193, 
        p_wishbone_n2194, p_wishbone_n2195, p_wishbone_n2196, p_wishbone_n2197, 
        p_wishbone_n2198, p_wishbone_n2199, p_wishbone_n2170, p_wishbone_n2201, 
        p_wishbone_n2202, p_wishbone_n2203, p_wishbone_n2204, p_wishbone_n2205, 
        p_wishbone_n2206, p_wishbone_n2207, p_wishbone_n2208, p_wishbone_n2209, 
        p_wishbone_n2210, p_wishbone_n2211, p_wishbone_n2212, p_wishbone_n2213, 
        p_wishbone_n2214, p_wishbone_n2215, p_wishbone_n2216, p_wishbone_n2217, 
        p_wishbone_n2218, p_wishbone_n2219, p_wishbone_n2220, p_wishbone_n2221, 
        p_wishbone_n2222, p_wishbone_n2223, p_wishbone_n2224, p_wishbone_n2225, 
        p_wishbone_n2226, p_wishbone_n2227, p_wishbone_n2228, p_wishbone_n2229, 
        p_wishbone_n2200, p_wishbone_n2339, p_wishbone_n2333, p_wishbone_n2334, 
        p_wishbone_n2342, p_wishbone_n2341, p_wishbone_n2335, p_wishbone_n2336, 
        p_wishbone_n2337, p_wishbone_n2340, p_wishbone_n2462, p_wishbone_n2250, 
        p_wishbone_n2258, p_wishbone_n2251, p_wishbone_n2259, p_wishbone_n2252, 
        p_wishbone_n2260, p_wishbone_n2253, p_wishbone_n2261, p_wishbone_n2254, 
        p_wishbone_n2262, p_wishbone_n2255, p_wishbone_n2263, p_wishbone_n2256, 
        p_wishbone_n2264, p_wishbone_n2257, p_wishbone_n2265, p_wishbone_n2266, 
        p_wishbone_n2267, p_wishbone_n2268, p_wishbone_n2269, p_wishbone_n2270, 
        p_wishbone_n2271, p_wishbone_n2272, p_wishbone_n2273, p_wishbone_n2274, 
        p_wishbone_n2275, p_wishbone_n2276, p_wishbone_n2277, p_wishbone_n2278, 
        p_wishbone_n2279, p_wishbone_n2280, p_wishbone_n2281, p_wishbone_n2282, 
        p_wishbone_n2283, p_wishbone_n2284, p_wishbone_n2285, p_wishbone_n2286, 
        p_wishbone_n2287, p_wishbone_n2288, p_wishbone_n2289, p_wishbone_n2290, 
        p_wishbone_n2291, p_wishbone_n2292, p_wishbone_n2293, 
        p_wishbone_TxStartFrm_syncb1, p_wishbone_TxStartFrm_sync2, 
        p_wishbone_TxStartFrm_sync1, p_wishbone_TxStartFrm_wb, 
        p_wishbone_n2294, p_wishbone_n2295, p_wishbone_n2437, p_wishbone_n2230, 
        p_wishbone_n2231, p_wishbone_n2249, n33933, 
        p_wishbone_BlockingTxStatusWrite_sync2, 
        p_wishbone_BlockingTxStatusWrite_sync1, 
        p_wishbone_BlockingTxStatusWrite, p_wishbone_n2232, p_wishbone_n2239, 
        p_wishbone_n2233, p_wishbone_n2241, p_wishbone_n2234, p_wishbone_n2242, 
        p_wishbone_n2235, p_wishbone_n2243, p_wishbone_n2236, p_wishbone_n2244, 
        p_wishbone_n2237, p_wishbone_n2245, p_wishbone_n2238, p_wishbone_n2246, 
        p_wishbone_n2247, p_wishbone_n2347, p_wishbone_n2240, p_wishbone_n2085, 
        p_wishbone_n2086, p_wishbone_n2441, p_wishbone_n2327, p_wishbone_n2328, 
        p_wishbone_n2329, p_wishbone_N75, p_wishbone_n2331, p_wishbone_n2469, 
        p_wishbone_n2456, p_wishbone_n2455, p_wishbone_n2454, p_wishbone_n2453, 
        p_wishbone_n2452, p_wishbone_n2451, p_wishbone_n2450, p_wishbone_n2449, 
        p_wishbone_n2448, p_wishbone_n2447, p_wishbone_n2446, p_wishbone_n2445, 
        p_wishbone_n2444, p_wishbone_n2443, p_wishbone_n2442, p_wishbone_n2440, 
        p_wishbone_n2439, p_wishbone_n2438, p_wishbone_n2436, p_wishbone_n2434, 
        p_wishbone_n2433, p_wishbone_n2432, p_wishbone_n2431, p_wishbone_n2430, 
        p_wishbone_n2429, p_wishbone_n2324, p_wishbone_n2323, p_wishbone_n2322, 
        p_wishbone_n2321, p_wishbone_n2087, p_wishbone_n2418, p_wishbone_n2419, 
        p_wishbone_n2420, p_wishbone_n2421, p_wishbone_n2422, p_wishbone_n2423, 
        p_wishbone_n2424, p_wishbone_n2088, p_wishbone_n2325, p_wishbone_n2382, 
        p_wishbone_n2406, p_wishbone_n2381, p_wishbone_n2405, p_wishbone_n2380, 
        p_wishbone_n2404, p_wishbone_n2379, p_wishbone_n2403, p_wishbone_n2378, 
        p_wishbone_n2402, p_wishbone_n2377, p_wishbone_n2401, p_wishbone_n2376, 
        p_wishbone_n2400, p_wishbone_n2375, p_wishbone_n2399, p_wishbone_n2365, 
        p_wishbone_n2366, p_wishbone_n2363, p_wishbone_n2364, p_wishbone_n2361, 
        p_wishbone_n2362, p_wishbone_n2359, p_wishbone_n2360, p_wishbone_n2357, 
        p_wishbone_n2358, p_wishbone_n2355, p_wishbone_n2356, p_wishbone_n2353, 
        p_wishbone_n2354, p_wishbone_n2351, p_wishbone_n2352, p_wishbone_n2373, 
        p_wishbone_n2372, p_wishbone_n2371, p_wishbone_n2370, p_wishbone_n2369, 
        p_wishbone_n2368, p_wishbone_n2367, p_wishbone_n2390, p_wishbone_n2389, 
        p_wishbone_n2388, p_wishbone_n2387, p_wishbone_n2386, p_wishbone_n2385, 
        p_wishbone_n2384, p_wishbone_n2383, p_wishbone_WriteRxDataToFifoSync2, 
        p_wishbone_WriteRxDataToFifoSync1, p_wishbone_WriteRxDataToFifo, 
        p_wishbone_n2413, p_wishbone_n2414, p_wishbone_n2411, p_wishbone_n2410, 
        p_wishbone_ShiftEndedSync_c1, p_wishbone_ShiftEndedSync2, 
        p_wishbone_ShiftEndedSync1, p_wishbone_ShiftEnded_rck, 
        p_wishbone_n2412, p_wishbone_n2407, p_wishbone_n2408, p_wishbone_n2409, 
        p_wishbone_n2425, p_wishbone_n2426, p_wishbone_n2427, p_wishbone_n2374, 
        p_wishbone_n2398, p_wishbone_n2397, p_wishbone_n2396, p_wishbone_n2395, 
        p_wishbone_n2394, p_wishbone_n2393, p_wishbone_n2392, p_wishbone_n2391, 
        p_wishbone_n2416, p_wishbone_n2415, p_wishbone_n2417, p_wishbone_n2326, 
        p_wishbone_RxEn, p_wishbone_n2428, p_wishbone_n2332, p_wishbone_WbEn, 
        p_wishbone_n2330, p_wishbone_n2089, p_wishbone_n2090, p_wishbone_n2091, 
        p_wishbone_n2092, p_wishbone_n2093, p_wishbone_n2094, p_wishbone_n2095, 
        p_wishbone_n2096, p_wishbone_n2097, p_wishbone_n2098, p_wishbone_n2099, 
        p_wishbone_n2100, p_wishbone_n2101, p_wishbone_n2102, p_wishbone_n2103, 
        p_wishbone_n2104, p_wishbone_n2248, p_wishbone_n2320, p_wishbone_n2301, 
        p_wishbone_n2302, p_wishbone_n2303, p_wishbone_n2304, p_wishbone_n2305, 
        p_wishbone_n2306, p_wishbone_n2307, p_wishbone_n2308, p_wishbone_n2309, 
        p_wishbone_n2310, p_wishbone_n2311, p_wishbone_n2312, p_wishbone_n2313, 
        p_wishbone_n2314, p_wishbone_n2299, p_wishbone_n2315, p_wishbone_n2316, 
        p_wishbone_n2105, p_wishbone_n2106, p_wishbone_n2107, p_wishbone_n2108, 
        p_wishbone_n2319, p_wishbone_TxEn, p_wishbone_n2457, p_wishbone_n2458, 
        p_wishbone_n2318, p_wishbone_n2317, p_wishbone_n2459, p_wishbone_n2460, 
        p_wishbone_n2461, p_wishbone_n2348, p_wishbone_N867, p_wishbone_n2349, 
        n33934, p_wishbone_n2463, p_wishbone_n2343, p_wishbone_n2344, 
        p_wishbone_n2345, p_wishbone_n2346, p_wishbone_n2350, p_wishbone_n2466, 
        p_wishbone_n2338, p_wishbone_n2464, p_wishbone_n2465, p_wishbone_n2467, 
        p_wishbone_ReadTxDataFromFifo_sync2, 
        p_wishbone_ReadTxDataFromFifo_syncb2, 
        p_wishbone_ReadTxDataFromFifo_syncb1, 
        p_wishbone_ReadTxDataFromFifo_sync1, p_wishbone_ReadTxDataFromFifo_tck, 
        p_wishbone_n2296, p_wishbone_n2297, p_wishbone_n2298, p_wishbone_n2300, 
        p_wishbone_LatchValidBytes, p_wishbone_N811, p_wishbone_n2468, 
        p_wishbone_n2435, p_wishbone_n2109, p_wishbone_n2470, p_wishbone_n2110, 
        p_wishbone_n2111, p_wishbone_n2112, p_wishbone_n2113, p_wishbone_n2114, 
        p_wishbone_n2115, p_wishbone_n2116, p_wishbone_n2117, p_wishbone_n2118, 
        p_wishbone_n2119, p_wishbone_n2120, p_wishbone_n2121, p_wishbone_n2122, 
        p_wishbone_n2123, p_wishbone_n2124, p_wishbone_n2125, p_wishbone_n2126, 
        p_wishbone_n2127, p_wishbone_n2128, p_wishbone_n2129, p_wishbone_n2130, 
        p_wishbone_n2131, p_wishbone_n2132, p_wishbone_n2133, 
        p_wishbone_RxAbortSyncb1, p_wishbone_RxAbortSync2, 
        p_wishbone_RxAbortSync3, p_wishbone_RxAbortSync1, 
        p_wishbone_RxAbortLatched, p_wishbone_n2471, p_wishbone_n2472, 
        p_wishbone_SyncRxStartFrm_q, p_wishbone_LatchedRxStartFrm, 
        p_wishbone_n2473, p_wishbone_TxAbort_wb, p_wishbone_TxAbortSync1, 
        TxAbort, p_wishbone_TxDone_wb, p_wishbone_TxDoneSync1, TxDone, 
        p_wishbone_TxRetry_wb, p_wishbone_TxRetrySync1, n33935, 
        p_wishbone_n2474, r_RxEn, r_TxEn, p_macstatus1_n89, p_macstatus1_n90, 
        p_macstatus1_n82, p_macstatus1_n83, p_macstatus1_n84, p_macstatus1_n85, 
        p_macstatus1_n86, p_macstatus1_n87, p_macstatus1_n91, p_macstatus1_n92, 
        p_macstatus1_n93, p_macstatus1_n94, p_macstatus1_n95, p_macstatus1_n96, 
        LoadRxStatus, p_macstatus1_TakeSample, p_macstatus1_N7, 
        p_macstatus1_n97, p_miim1_clkgen_n35, p_miim1_clkgen_N21, 
        p_miim1_clkgen_N20, p_miim1_clkgen_N19, p_miim1_clkgen_N18, 
        p_miim1_clkgen_N17, p_miim1_clkgen_N16, p_miim1_clkgen_N15, 
        p_miim1_shftrg_n145, p_miim1_shftrg_n146, p_miim1_shftrg_n147, 
        p_miim1_shftrg_n148, p_miim1_shftrg_n149, p_miim1_shftrg_n150, 
        p_miim1_shftrg_n151, p_miim1_shftrg_n152, p_miim1_shftrg_n153, 
        p_miim1_shftrg_n154, p_miim1_shftrg_n155, p_miim1_shftrg_n156, 
        p_miim1_shftrg_n157, p_miim1_shftrg_n158, p_miim1_shftrg_n159, 
        p_miim1_shftrg_n160, p_miim1_shftrg_n161, p_miim1_shftrg_n137, 
        p_miim1_shftrg_n138, p_miim1_shftrg_n139, p_miim1_shftrg_n140, 
        p_miim1_shftrg_n141, p_miim1_shftrg_n142, p_miim1_shftrg_n143, 
        p_miim1_shftrg_n144, p_miim1_outctrl_n33, p_miim1_outctrl_n34, 
        p_miim1_outctrl_n35, p_miim1_outctrl_n36, p_miim1_outctrl_n37, 
        p_miim1_outctrl_n38, p_ethreg1_MODER_0_n21, p_ethreg1_MODER_0_n22, 
        p_ethreg1_MODER_0_n23, p_ethreg1_MODER_0_n24, p_ethreg1_MODER_0_n25, 
        p_ethreg1_MODER_0_n26, p_ethreg1_MODER_0_n27, p_ethreg1_MODER_0_n28, 
        p_ethreg1_MODER_1_n23, p_ethreg1_MODER_1_n24, p_ethreg1_MODER_1_n25, 
        p_ethreg1_MODER_1_n26, p_ethreg1_MODER_1_n27, n33922, 
        p_ethreg1_MODER_1_n29, n33921, n33920, p_ethreg1_INT_MASK_0_n19, 
        p_ethreg1_INT_MASK_0_n20, p_ethreg1_INT_MASK_0_n21, 
        p_ethreg1_INT_MASK_0_n22, p_ethreg1_INT_MASK_0_n23, 
        p_ethreg1_INT_MASK_0_n24, p_ethreg1_INT_MASK_0_n25, 
        p_ethreg1_IPGT_0_n21, n33931, p_ethreg1_IPGT_0_n23, 
        p_ethreg1_IPGT_0_n24, n33927, p_ethreg1_IPGT_0_n26, 
        p_ethreg1_IPGT_0_n27, p_ethreg1_IPGR1_0_n21, p_ethreg1_IPGR1_0_n22, 
        n33929, n33928, p_ethreg1_IPGR1_0_n25, p_ethreg1_IPGR1_0_n26, 
        p_ethreg1_IPGR1_0_n27, p_ethreg1_PACKETLEN_1_n23, n33924, n33923, 
        p_ethreg1_PACKETLEN_1_n26, p_ethreg1_PACKETLEN_1_n27, 
        p_ethreg1_PACKETLEN_1_n28, p_ethreg1_PACKETLEN_1_n29, 
        p_ethreg1_PACKETLEN_1_n30, p_ethreg1_PACKETLEN_2_n22, 
        p_ethreg1_PACKETLEN_2_n23, p_ethreg1_PACKETLEN_2_n24, 
        p_ethreg1_PACKETLEN_2_n25, p_ethreg1_PACKETLEN_2_n26, 
        p_ethreg1_PACKETLEN_2_n27, p_ethreg1_PACKETLEN_2_n17, 
        p_ethreg1_PACKETLEN_2_n29, p_ethreg1_COLLCONF_0_n21, 
        p_ethreg1_COLLCONF_0_n22, p_ethreg1_COLLCONF_0_n23, 
        p_ethreg1_COLLCONF_0_n24, p_ethreg1_COLLCONF_0_n25, 
        p_ethreg1_COLLCONF_0_n26, p_ethreg1_COLLCONF_2_n15, 
        p_ethreg1_COLLCONF_2_n16, p_ethreg1_COLLCONF_2_n17, 
        p_ethreg1_COLLCONF_2_n18, p_ethreg1_CTRLMODER_0_n10, 
        p_ethreg1_CTRLMODER_0_n11, p_ethreg1_CTRLMODER_0_n12, 
        p_ethreg1_MIIMODER_0_n24, p_ethreg1_MIIMODER_0_n25, 
        p_ethreg1_MIIMODER_0_n26, p_ethreg1_MIIMODER_0_n27, 
        p_ethreg1_MIIMODER_0_n28, p_ethreg1_MIIMODER_0_n29, 
        p_ethreg1_MIIMODER_0_n30, p_ethreg1_MIIMODER_0_n31, n33932, 
        p_ethreg1_MIIADDRESS_0_n15, p_ethreg1_MIIADDRESS_0_n16, 
        p_ethreg1_MIIADDRESS_0_n17, p_ethreg1_MIIADDRESS_0_n18, 
        p_ethreg1_MIIADDRESS_0_n19, p_ethreg1_MIIRX_DATA_n37, 
        p_ethreg1_MIIRX_DATA_n38, p_ethreg1_MIIRX_DATA_n39, 
        p_ethreg1_MIIRX_DATA_n40, p_ethreg1_MIIRX_DATA_n41, 
        p_ethreg1_MIIRX_DATA_n42, p_ethreg1_MIIRX_DATA_n43, 
        p_ethreg1_MIIRX_DATA_n44, p_ethreg1_MIIRX_DATA_n45, 
        p_ethreg1_MIIRX_DATA_n46, p_ethreg1_MIIRX_DATA_n47, 
        p_ethreg1_MIIRX_DATA_n48, p_ethreg1_MIIRX_DATA_n49, 
        p_ethreg1_MIIRX_DATA_n50, p_ethreg1_MIIRX_DATA_n51, 
        p_ethreg1_MIIRX_DATA_n52, p_maccontrol1_receivecontrol1_n503, 
        p_maccontrol1_receivecontrol1_n507, p_maccontrol1_receivecontrol1_n506, 
        p_maccontrol1_receivecontrol1_n505, p_maccontrol1_receivecontrol1_n504, 
        p_maccontrol1_receivecontrol1_n524, p_maccontrol1_receivecontrol1_n501, 
        p_maccontrol1_receivecontrol1_PauseTimerEq0_sync1, n33939, 
        p_maccontrol1_receivecontrol1_N208, p_maccontrol1_receivecontrol1_n508, 
        p_maccontrol1_receivecontrol1_n509, p_maccontrol1_receivecontrol1_n510, 
        p_maccontrol1_receivecontrol1_n511, p_maccontrol1_receivecontrol1_n512, 
        p_maccontrol1_receivecontrol1_n513, p_maccontrol1_receivecontrol1_n514, 
        p_maccontrol1_receivecontrol1_n515, p_maccontrol1_receivecontrol1_n516, 
        p_maccontrol1_receivecontrol1_n517, p_maccontrol1_receivecontrol1_n518, 
        p_maccontrol1_receivecontrol1_n519, p_maccontrol1_receivecontrol1_n520, 
        p_maccontrol1_receivecontrol1_n521, p_maccontrol1_receivecontrol1_n522, 
        p_maccontrol1_receivecontrol1_n523, p_maccontrol1_receivecontrol1_n525, 
        p_maccontrol1_receivecontrol1_n541, p_maccontrol1_receivecontrol1_n540, 
        p_maccontrol1_receivecontrol1_n539, p_maccontrol1_receivecontrol1_n538, 
        p_maccontrol1_receivecontrol1_n537, p_maccontrol1_receivecontrol1_n536, 
        p_maccontrol1_receivecontrol1_n535, p_maccontrol1_receivecontrol1_n534, 
        p_maccontrol1_receivecontrol1_n533, p_maccontrol1_receivecontrol1_n532, 
        p_maccontrol1_receivecontrol1_n531, p_maccontrol1_receivecontrol1_n530, 
        p_maccontrol1_receivecontrol1_n529, p_maccontrol1_receivecontrol1_n528, 
        p_maccontrol1_receivecontrol1_n527, p_maccontrol1_receivecontrol1_n526, 
        p_maccontrol1_receivecontrol1_n558, p_maccontrol1_receivecontrol1_n559, 
        p_maccontrol1_receivecontrol1_n561, p_maccontrol1_receivecontrol1_n560, 
        p_maccontrol1_receivecontrol1_n557, p_maccontrol1_receivecontrol1_n556, 
        p_maccontrol1_receivecontrol1_n555, p_maccontrol1_receivecontrol1_n554, 
        p_maccontrol1_receivecontrol1_n553, p_maccontrol1_receivecontrol1_n552, 
        p_maccontrol1_receivecontrol1_n551, p_maccontrol1_receivecontrol1_n550, 
        p_maccontrol1_receivecontrol1_n549, p_maccontrol1_receivecontrol1_n548, 
        p_maccontrol1_receivecontrol1_n547, p_maccontrol1_receivecontrol1_n546, 
        p_maccontrol1_receivecontrol1_n545, p_maccontrol1_receivecontrol1_n544, 
        p_maccontrol1_receivecontrol1_n543, p_maccontrol1_receivecontrol1_n542, 
        p_maccontrol1_receivecontrol1_n564, p_maccontrol1_receivecontrol1_n563, 
        p_maccontrol1_receivecontrol1_n562, p_maccontrol1_receivecontrol1_n566, 
        p_maccontrol1_receivecontrol1_n565, p_maccontrol1_receivecontrol1_n567, 
        p_maccontrol1_receivecontrol1_n568, p_maccontrol1_receivecontrol1_n569, 
        p_maccontrol1_receivecontrol1_n570, 
        p_maccontrol1_transmitcontrol1_n263, 
        p_maccontrol1_transmitcontrol1_n264, 
        p_maccontrol1_transmitcontrol1_n265, 
        p_maccontrol1_transmitcontrol1_n266, 
        p_maccontrol1_transmitcontrol1_n267, 
        p_maccontrol1_transmitcontrol1_n268, 
        p_maccontrol1_transmitcontrol1_n269, 
        p_maccontrol1_transmitcontrol1_n270, 
        p_maccontrol1_transmitcontrol1_n275, 
        p_maccontrol1_transmitcontrol1_n274, 
        p_maccontrol1_transmitcontrol1_n273, 
        p_maccontrol1_transmitcontrol1_n272, 
        p_maccontrol1_transmitcontrol1_n283, 
        p_maccontrol1_transmitcontrol1_n276, 
        p_maccontrol1_transmitcontrol1_n277, 
        p_maccontrol1_transmitcontrol1_n278, 
        p_maccontrol1_transmitcontrol1_n279, 
        p_maccontrol1_transmitcontrol1_n271, p_maccontrol1_TxCtrlStartFrm, 
        p_maccontrol1_transmitcontrol1_n280, 
        p_maccontrol1_transmitcontrol1_n281, 
        p_maccontrol1_transmitcontrol1_n282, 
        p_maccontrol1_transmitcontrol1_N31, 
        p_maccontrol1_transmitcontrol1_n285, 
        p_maccontrol1_transmitcontrol1_n284, p_txethmac1_txcounters1_n172, 
        p_txethmac1_txcounters1_n173, p_txethmac1_txcounters1_n174, 
        p_txethmac1_txcounters1_n188, p_txethmac1_txcounters1_n187, 
        p_txethmac1_txcounters1_n186, p_txethmac1_txcounters1_n185, 
        p_txethmac1_txcounters1_n184, p_txethmac1_txcounters1_n183, 
        p_txethmac1_txcounters1_n182, p_txethmac1_txcounters1_n181, 
        p_txethmac1_txcounters1_n180, p_txethmac1_txcounters1_n179, 
        p_txethmac1_txcounters1_n178, p_txethmac1_txcounters1_n177, 
        p_txethmac1_txcounters1_n176, p_txethmac1_txcounters1_n175, 
        p_txethmac1_txcounters1_n189, p_txethmac1_txcounters1_n190, 
        p_txethmac1_txcounters1_n191, p_txethmac1_txcounters1_n192, 
        p_txethmac1_txcounters1_n193, p_txethmac1_txcounters1_n194, 
        p_txethmac1_txcounters1_n195, p_txethmac1_txcounters1_n196, 
        p_txethmac1_txcounters1_n197, p_txethmac1_txcounters1_n198, 
        p_txethmac1_txcounters1_n199, p_txethmac1_txcounters1_n200, 
        p_txethmac1_txcounters1_n201, p_txethmac1_txcounters1_n202, 
        p_txethmac1_txcounters1_n204, p_txethmac1_txcounters1_n203, 
        p_txethmac1_txcounters1_n205, p_txethmac1_txcounters1_n206, 
        p_txethmac1_txstatem1_n90, p_txethmac1_StateJam, 
        p_txethmac1_txstatem1_n93, p_txethmac1_txstatem1_n94, 
        p_txethmac1_StartData_1, p_txethmac1_StartData_0, 
        p_txethmac1_txstatem1_n95, p_txethmac1_txstatem1_n96, 
        p_txethmac1_txstatem1_n97, p_txethmac1_txstatem1_n92, 
        p_txethmac1_txstatem1_n91, p_txethmac1_txstatem1_n98, 
        p_txethmac1_txcrc_N25, p_txethmac1_txcrc_N21, p_txethmac1_txcrc_N17, 
        p_txethmac1_txcrc_N13, p_txethmac1_txcrc_N9, p_txethmac1_txcrc_N5, 
        p_txethmac1_txcrc_N8, p_txethmac1_txcrc_N26, p_txethmac1_txcrc_N22, 
        p_txethmac1_txcrc_N18, p_txethmac1_txcrc_N14, p_txethmac1_txcrc_N10, 
        p_txethmac1_txcrc_N6, p_txethmac1_txcrc_N34, p_txethmac1_txcrc_N30, 
        p_txethmac1_txcrc_N4, p_txethmac1_txcrc_N32, p_txethmac1_txcrc_N28, 
        p_txethmac1_txcrc_N24, p_txethmac1_txcrc_N20, p_txethmac1_txcrc_N16, 
        p_txethmac1_txcrc_N12, p_txethmac1_txcrc_N33, p_txethmac1_txcrc_N29, 
        p_txethmac1_txcrc_N31, p_txethmac1_txcrc_N27, p_txethmac1_txcrc_N23, 
        p_txethmac1_txcrc_N19, p_txethmac1_txcrc_N15, p_txethmac1_txcrc_N11, 
        p_txethmac1_txcrc_N7, p_txethmac1_txcrc_N3, p_txethmac1_random1_n98, 
        p_txethmac1_random1_n99, p_txethmac1_random1_n100, 
        p_txethmac1_random1_n101, p_txethmac1_random1_n102, 
        p_txethmac1_random1_n103, p_txethmac1_random1_n104, 
        p_txethmac1_random1_n105, p_txethmac1_random1_n106, 
        p_txethmac1_random1_n107, p_txethmac1_random1_x_8, 
        p_txethmac1_random1_x_7, p_txethmac1_random1_x_6, 
        p_txethmac1_random1_x_5, p_txethmac1_random1_x_4, 
        p_txethmac1_random1_x_3, p_txethmac1_random1_x_2, 
        p_txethmac1_random1_x_1, p_txethmac1_random1_x_0, 
        p_txethmac1_random1_n108, p_rxethmac1_rxstatem1_n38, 
        p_rxethmac1_rxstatem1_n37, p_rxethmac1_rxstatem1_n39, 
        p_rxethmac1_rxstatem1_n40, p_rxethmac1_rxstatem1_n41, 
        p_rxethmac1_rxstatem1_n42, p_rxethmac1_rxcounters1_n175, 
        p_rxethmac1_rxcounters1_n174, p_rxethmac1_rxcounters1_n173, 
        p_rxethmac1_rxcounters1_n172, p_rxethmac1_rxcounters1_n171, 
        p_rxethmac1_rxcounters1_n170, p_rxethmac1_rxcounters1_n169, 
        p_rxethmac1_rxcounters1_n168, p_rxethmac1_rxcounters1_n167, 
        p_rxethmac1_rxcounters1_n166, p_rxethmac1_rxcounters1_n165, 
        p_rxethmac1_rxcounters1_n164, p_rxethmac1_rxcounters1_n163, 
        p_rxethmac1_rxcounters1_n162, p_rxethmac1_rxcounters1_n176, 
        p_rxethmac1_rxcounters1_n161, p_rxethmac1_rxcounters1_n178, 
        p_rxethmac1_rxcounters1_n177, p_rxethmac1_rxcounters1_n179, 
        p_rxethmac1_rxcounters1_n180, p_rxethmac1_rxcounters1_n183, 
        p_rxethmac1_rxcounters1_n182, p_rxethmac1_rxcounters1_n181, 
        p_rxethmac1_rxcounters1_n184, p_rxethmac1_rxcounters1_n185, 
        p_rxethmac1_rxaddrcheck1_n290, p_rxethmac1_rxaddrcheck1_n294, 
        p_rxethmac1_rxaddrcheck1_N10, p_rxethmac1_rxaddrcheck1_n295, 
        p_wishbone_bd_ram_n17793, p_wishbone_bd_ram_n17794, 
        p_wishbone_bd_ram_n17795, p_wishbone_bd_ram_n17796, 
        p_wishbone_bd_ram_n17797, p_wishbone_bd_ram_n17798, 
        p_wishbone_bd_ram_n17799, p_wishbone_bd_ram_n17800, 
        p_wishbone_bd_ram_n17801, p_wishbone_bd_ram_n17802, 
        p_wishbone_bd_ram_n17803, p_wishbone_bd_ram_n17804, 
        p_wishbone_bd_ram_n17805, p_wishbone_bd_ram_n17806, 
        p_wishbone_bd_ram_n17807, p_wishbone_bd_ram_n17808, 
        p_wishbone_bd_ram_n17809, p_wishbone_bd_ram_n17810, 
        p_wishbone_bd_ram_n17811, p_wishbone_bd_ram_n17812, 
        p_wishbone_bd_ram_n17813, p_wishbone_bd_ram_n17814, 
        p_wishbone_bd_ram_n17815, p_wishbone_bd_ram_n17816, 
        p_wishbone_bd_ram_n17817, p_wishbone_bd_ram_n17818, 
        p_wishbone_bd_ram_n17819, p_wishbone_bd_ram_n17820, 
        p_wishbone_bd_ram_n17821, p_wishbone_bd_ram_n17822, 
        p_wishbone_bd_ram_n17823, p_wishbone_bd_ram_n17824, 
        p_wishbone_bd_ram_n17825, p_wishbone_bd_ram_n17826, 
        p_wishbone_bd_ram_n17827, p_wishbone_bd_ram_n17828, 
        p_wishbone_bd_ram_n17829, p_wishbone_bd_ram_n17830, 
        p_wishbone_bd_ram_n17831, p_wishbone_bd_ram_n17832, 
        p_wishbone_bd_ram_n17833, p_wishbone_bd_ram_n17834, 
        p_wishbone_bd_ram_n17835, p_wishbone_bd_ram_n17836, 
        p_wishbone_bd_ram_n17837, p_wishbone_bd_ram_n17838, 
        p_wishbone_bd_ram_n17839, p_wishbone_bd_ram_n17840, 
        p_wishbone_bd_ram_n17841, p_wishbone_bd_ram_n17842, 
        p_wishbone_bd_ram_n17843, p_wishbone_bd_ram_n17844, 
        p_wishbone_bd_ram_n17845, p_wishbone_bd_ram_n17846, 
        p_wishbone_bd_ram_n17847, p_wishbone_bd_ram_n17848, 
        p_wishbone_bd_ram_n17849, p_wishbone_bd_ram_n17850, 
        p_wishbone_bd_ram_n17851, p_wishbone_bd_ram_n17852, 
        p_wishbone_bd_ram_n17853, p_wishbone_bd_ram_n17854, 
        p_wishbone_bd_ram_n17855, p_wishbone_bd_ram_n17856, 
        p_wishbone_bd_ram_n17857, p_wishbone_bd_ram_n17858, 
        p_wishbone_bd_ram_n17859, p_wishbone_bd_ram_n17860, 
        p_wishbone_bd_ram_n17861, p_wishbone_bd_ram_n17862, 
        p_wishbone_bd_ram_n17863, p_wishbone_bd_ram_n17864, 
        p_wishbone_bd_ram_n17865, p_wishbone_bd_ram_n17866, 
        p_wishbone_bd_ram_n17867, p_wishbone_bd_ram_n17868, 
        p_wishbone_bd_ram_n17869, p_wishbone_bd_ram_n17870, 
        p_wishbone_bd_ram_n17871, p_wishbone_bd_ram_n17872, 
        p_wishbone_bd_ram_n17873, p_wishbone_bd_ram_n17874, 
        p_wishbone_bd_ram_n17875, p_wishbone_bd_ram_n17876, 
        p_wishbone_bd_ram_n17877, p_wishbone_bd_ram_n17878, 
        p_wishbone_bd_ram_n17879, p_wishbone_bd_ram_n17880, 
        p_wishbone_bd_ram_n17881, p_wishbone_bd_ram_n17882, 
        p_wishbone_bd_ram_n17883, p_wishbone_bd_ram_n17884, 
        p_wishbone_bd_ram_n17885, p_wishbone_bd_ram_n17886, 
        p_wishbone_bd_ram_n17887, p_wishbone_bd_ram_n17888, 
        p_wishbone_bd_ram_n17889, p_wishbone_bd_ram_n17890, 
        p_wishbone_bd_ram_n17891, p_wishbone_bd_ram_n17892, 
        p_wishbone_bd_ram_n17893, p_wishbone_bd_ram_n17894, 
        p_wishbone_bd_ram_n17895, p_wishbone_bd_ram_n17896, 
        p_wishbone_bd_ram_n17897, p_wishbone_bd_ram_n17898, 
        p_wishbone_bd_ram_n17899, p_wishbone_bd_ram_n17900, 
        p_wishbone_bd_ram_n17901, p_wishbone_bd_ram_n17902, 
        p_wishbone_bd_ram_n17903, p_wishbone_bd_ram_n17904, 
        p_wishbone_bd_ram_n17905, p_wishbone_bd_ram_n17906, 
        p_wishbone_bd_ram_n17907, p_wishbone_bd_ram_n17908, 
        p_wishbone_bd_ram_n17909, p_wishbone_bd_ram_n17910, 
        p_wishbone_bd_ram_n17911, p_wishbone_bd_ram_n17912, 
        p_wishbone_bd_ram_n17913, p_wishbone_bd_ram_n17914, 
        p_wishbone_bd_ram_n17915, p_wishbone_bd_ram_n17916, 
        p_wishbone_bd_ram_n17917, p_wishbone_bd_ram_n17918, 
        p_wishbone_bd_ram_n17919, p_wishbone_bd_ram_n17920, 
        p_wishbone_bd_ram_n17921, p_wishbone_bd_ram_n17922, 
        p_wishbone_bd_ram_n17923, p_wishbone_bd_ram_n17924, 
        p_wishbone_bd_ram_n17925, p_wishbone_bd_ram_n17926, 
        p_wishbone_bd_ram_n17927, p_wishbone_bd_ram_n17928, 
        p_wishbone_bd_ram_n17929, p_wishbone_bd_ram_n17930, 
        p_wishbone_bd_ram_n17931, p_wishbone_bd_ram_n17932, 
        p_wishbone_bd_ram_n17933, p_wishbone_bd_ram_n17934, 
        p_wishbone_bd_ram_n17935, p_wishbone_bd_ram_n17936, 
        p_wishbone_bd_ram_n17937, p_wishbone_bd_ram_n17938, 
        p_wishbone_bd_ram_n17939, p_wishbone_bd_ram_n17940, 
        p_wishbone_bd_ram_n17941, p_wishbone_bd_ram_n17942, 
        p_wishbone_bd_ram_n17943, p_wishbone_bd_ram_n17944, 
        p_wishbone_bd_ram_n17945, p_wishbone_bd_ram_n17946, 
        p_wishbone_bd_ram_n17947, p_wishbone_bd_ram_n17948, 
        p_wishbone_bd_ram_n17949, p_wishbone_bd_ram_n17950, 
        p_wishbone_bd_ram_n17951, p_wishbone_bd_ram_n17952, 
        p_wishbone_bd_ram_n17953, p_wishbone_bd_ram_n17954, 
        p_wishbone_bd_ram_n17955, p_wishbone_bd_ram_n17956, 
        p_wishbone_bd_ram_n17957, p_wishbone_bd_ram_n17958, 
        p_wishbone_bd_ram_n17959, p_wishbone_bd_ram_n17960, 
        p_wishbone_bd_ram_n17961, p_wishbone_bd_ram_n17962, 
        p_wishbone_bd_ram_n17963, p_wishbone_bd_ram_n17964, 
        p_wishbone_bd_ram_n17965, p_wishbone_bd_ram_n17966, 
        p_wishbone_bd_ram_n17967, p_wishbone_bd_ram_n17968, 
        p_wishbone_bd_ram_n17969, p_wishbone_bd_ram_n17970, 
        p_wishbone_bd_ram_n17971, p_wishbone_bd_ram_n17972, 
        p_wishbone_bd_ram_n17973, p_wishbone_bd_ram_n17974, 
        p_wishbone_bd_ram_n17975, p_wishbone_bd_ram_n17976, 
        p_wishbone_bd_ram_n17977, p_wishbone_bd_ram_n17978, 
        p_wishbone_bd_ram_n17979, p_wishbone_bd_ram_n17980, 
        p_wishbone_bd_ram_n17981, p_wishbone_bd_ram_n17982, 
        p_wishbone_bd_ram_n17983, p_wishbone_bd_ram_n17984, 
        p_wishbone_bd_ram_n17985, p_wishbone_bd_ram_n17986, 
        p_wishbone_bd_ram_n17987, p_wishbone_bd_ram_n17988, 
        p_wishbone_bd_ram_n17989, p_wishbone_bd_ram_n17990, 
        p_wishbone_bd_ram_n17991, p_wishbone_bd_ram_n17992, 
        p_wishbone_bd_ram_n17993, p_wishbone_bd_ram_n17994, 
        p_wishbone_bd_ram_n17995, p_wishbone_bd_ram_n17996, 
        p_wishbone_bd_ram_n17997, p_wishbone_bd_ram_n17998, 
        p_wishbone_bd_ram_n17999, p_wishbone_bd_ram_n18000, 
        p_wishbone_bd_ram_n18001, p_wishbone_bd_ram_n18002, 
        p_wishbone_bd_ram_n18003, p_wishbone_bd_ram_n18004, 
        p_wishbone_bd_ram_n18005, p_wishbone_bd_ram_n18006, 
        p_wishbone_bd_ram_n18007, p_wishbone_bd_ram_n18008, 
        p_wishbone_bd_ram_n18009, p_wishbone_bd_ram_n18010, 
        p_wishbone_bd_ram_n18011, p_wishbone_bd_ram_n18012, 
        p_wishbone_bd_ram_n18013, p_wishbone_bd_ram_n18014, 
        p_wishbone_bd_ram_n18015, p_wishbone_bd_ram_n18016, 
        p_wishbone_bd_ram_n18017, p_wishbone_bd_ram_n18018, 
        p_wishbone_bd_ram_n18019, p_wishbone_bd_ram_n18020, 
        p_wishbone_bd_ram_n18021, p_wishbone_bd_ram_n18022, 
        p_wishbone_bd_ram_n18023, p_wishbone_bd_ram_n18024, 
        p_wishbone_bd_ram_n18025, p_wishbone_bd_ram_n18026, 
        p_wishbone_bd_ram_n18027, p_wishbone_bd_ram_n18028, 
        p_wishbone_bd_ram_n18029, p_wishbone_bd_ram_n18030, 
        p_wishbone_bd_ram_n18031, p_wishbone_bd_ram_n18032, 
        p_wishbone_bd_ram_n18033, p_wishbone_bd_ram_n18034, 
        p_wishbone_bd_ram_n18035, p_wishbone_bd_ram_n18036, 
        p_wishbone_bd_ram_n18037, p_wishbone_bd_ram_n18038, 
        p_wishbone_bd_ram_n18039, p_wishbone_bd_ram_n18040, 
        p_wishbone_bd_ram_n18041, p_wishbone_bd_ram_n18042, 
        p_wishbone_bd_ram_n18043, p_wishbone_bd_ram_n18044, 
        p_wishbone_bd_ram_n18045, p_wishbone_bd_ram_n18046, 
        p_wishbone_bd_ram_n18047, p_wishbone_bd_ram_n18048, 
        p_wishbone_bd_ram_n18049, p_wishbone_bd_ram_n18050, 
        p_wishbone_bd_ram_n18051, p_wishbone_bd_ram_n18052, 
        p_wishbone_bd_ram_n18053, p_wishbone_bd_ram_n18054, 
        p_wishbone_bd_ram_n18055, p_wishbone_bd_ram_n18056, 
        p_wishbone_bd_ram_n18057, p_wishbone_bd_ram_n18058, 
        p_wishbone_bd_ram_n18059, p_wishbone_bd_ram_n18060, 
        p_wishbone_bd_ram_n18061, p_wishbone_bd_ram_n18062, 
        p_wishbone_bd_ram_n18063, p_wishbone_bd_ram_n18064, 
        p_wishbone_bd_ram_n18065, p_wishbone_bd_ram_n18066, 
        p_wishbone_bd_ram_n18067, p_wishbone_bd_ram_n18068, 
        p_wishbone_bd_ram_n18069, p_wishbone_bd_ram_n18070, 
        p_wishbone_bd_ram_n18071, p_wishbone_bd_ram_n18072, 
        p_wishbone_bd_ram_n18073, p_wishbone_bd_ram_n18074, 
        p_wishbone_bd_ram_n18075, p_wishbone_bd_ram_n18076, 
        p_wishbone_bd_ram_n18077, p_wishbone_bd_ram_n18078, 
        p_wishbone_bd_ram_n18079, p_wishbone_bd_ram_n18080, 
        p_wishbone_bd_ram_n18081, p_wishbone_bd_ram_n18082, 
        p_wishbone_bd_ram_n18083, p_wishbone_bd_ram_n18084, 
        p_wishbone_bd_ram_n18085, p_wishbone_bd_ram_n18086, 
        p_wishbone_bd_ram_n18087, p_wishbone_bd_ram_n18088, 
        p_wishbone_bd_ram_n18089, p_wishbone_bd_ram_n18090, 
        p_wishbone_bd_ram_n18091, p_wishbone_bd_ram_n18092, 
        p_wishbone_bd_ram_n18093, p_wishbone_bd_ram_n18094, 
        p_wishbone_bd_ram_n18095, p_wishbone_bd_ram_n18096, 
        p_wishbone_bd_ram_n18097, p_wishbone_bd_ram_n18098, 
        p_wishbone_bd_ram_n18099, p_wishbone_bd_ram_n18100, 
        p_wishbone_bd_ram_n18101, p_wishbone_bd_ram_n18102, 
        p_wishbone_bd_ram_n18103, p_wishbone_bd_ram_n18104, 
        p_wishbone_bd_ram_n18105, p_wishbone_bd_ram_n18106, 
        p_wishbone_bd_ram_n18107, p_wishbone_bd_ram_n18108, 
        p_wishbone_bd_ram_n18109, p_wishbone_bd_ram_n18110, 
        p_wishbone_bd_ram_n18111, p_wishbone_bd_ram_n18112, 
        p_wishbone_bd_ram_n18113, p_wishbone_bd_ram_n18114, 
        p_wishbone_bd_ram_n18115, p_wishbone_bd_ram_n18116, 
        p_wishbone_bd_ram_n18117, p_wishbone_bd_ram_n18118, 
        p_wishbone_bd_ram_n18119, p_wishbone_bd_ram_n18120, 
        p_wishbone_bd_ram_n18121, p_wishbone_bd_ram_n18122, 
        p_wishbone_bd_ram_n18123, p_wishbone_bd_ram_n18124, 
        p_wishbone_bd_ram_n18125, p_wishbone_bd_ram_n18126, 
        p_wishbone_bd_ram_n18127, p_wishbone_bd_ram_n18128, 
        p_wishbone_bd_ram_n18129, p_wishbone_bd_ram_n18130, 
        p_wishbone_bd_ram_n18131, p_wishbone_bd_ram_n18132, 
        p_wishbone_bd_ram_n18133, p_wishbone_bd_ram_n18134, 
        p_wishbone_bd_ram_n18135, p_wishbone_bd_ram_n18136, 
        p_wishbone_bd_ram_n18137, p_wishbone_bd_ram_n18138, 
        p_wishbone_bd_ram_n18139, p_wishbone_bd_ram_n18140, 
        p_wishbone_bd_ram_n18141, p_wishbone_bd_ram_n18142, 
        p_wishbone_bd_ram_n18143, p_wishbone_bd_ram_n18144, 
        p_wishbone_bd_ram_n18145, p_wishbone_bd_ram_n18146, 
        p_wishbone_bd_ram_n18147, p_wishbone_bd_ram_n18148, 
        p_wishbone_bd_ram_n18149, p_wishbone_bd_ram_n18150, 
        p_wishbone_bd_ram_n18151, p_wishbone_bd_ram_n18152, 
        p_wishbone_bd_ram_n18153, p_wishbone_bd_ram_n18154, 
        p_wishbone_bd_ram_n18155, p_wishbone_bd_ram_n18156, 
        p_wishbone_bd_ram_n18157, p_wishbone_bd_ram_n18158, 
        p_wishbone_bd_ram_n18159, p_wishbone_bd_ram_n18160, 
        p_wishbone_bd_ram_n18161, p_wishbone_bd_ram_n18162, 
        p_wishbone_bd_ram_n18163, p_wishbone_bd_ram_n18164, 
        p_wishbone_bd_ram_n18165, p_wishbone_bd_ram_n18166, 
        p_wishbone_bd_ram_n18167, p_wishbone_bd_ram_n18168, 
        p_wishbone_bd_ram_n18169, p_wishbone_bd_ram_n18170, 
        p_wishbone_bd_ram_n18171, p_wishbone_bd_ram_n18172, 
        p_wishbone_bd_ram_n18173, p_wishbone_bd_ram_n18174, 
        p_wishbone_bd_ram_n18175, p_wishbone_bd_ram_n18176, 
        p_wishbone_bd_ram_n18177, p_wishbone_bd_ram_n18178, 
        p_wishbone_bd_ram_n18179, p_wishbone_bd_ram_n18180, 
        p_wishbone_bd_ram_n18181, p_wishbone_bd_ram_n18182, 
        p_wishbone_bd_ram_n18183, p_wishbone_bd_ram_n18184, 
        p_wishbone_bd_ram_n18185, p_wishbone_bd_ram_n18186, 
        p_wishbone_bd_ram_n18187, p_wishbone_bd_ram_n18188, 
        p_wishbone_bd_ram_n18189, p_wishbone_bd_ram_n18190, 
        p_wishbone_bd_ram_n18191, p_wishbone_bd_ram_n18192, 
        p_wishbone_bd_ram_n18193, p_wishbone_bd_ram_n18194, 
        p_wishbone_bd_ram_n18195, p_wishbone_bd_ram_n18196, 
        p_wishbone_bd_ram_n18197, p_wishbone_bd_ram_n18198, 
        p_wishbone_bd_ram_n18199, p_wishbone_bd_ram_n18200, 
        p_wishbone_bd_ram_n18201, p_wishbone_bd_ram_n18202, 
        p_wishbone_bd_ram_n18203, p_wishbone_bd_ram_n18204, 
        p_wishbone_bd_ram_n18205, p_wishbone_bd_ram_n18206, 
        p_wishbone_bd_ram_n18207, p_wishbone_bd_ram_n18208, 
        p_wishbone_bd_ram_n18209, p_wishbone_bd_ram_n18210, 
        p_wishbone_bd_ram_n18211, p_wishbone_bd_ram_n18212, 
        p_wishbone_bd_ram_n18213, p_wishbone_bd_ram_n18214, 
        p_wishbone_bd_ram_n18215, p_wishbone_bd_ram_n18216, 
        p_wishbone_bd_ram_n18217, p_wishbone_bd_ram_n18218, 
        p_wishbone_bd_ram_n18219, p_wishbone_bd_ram_n18220, 
        p_wishbone_bd_ram_n18221, p_wishbone_bd_ram_n18222, 
        p_wishbone_bd_ram_n18223, p_wishbone_bd_ram_n18224, 
        p_wishbone_bd_ram_n18225, p_wishbone_bd_ram_n18226, 
        p_wishbone_bd_ram_n18227, p_wishbone_bd_ram_n18228, 
        p_wishbone_bd_ram_n18229, p_wishbone_bd_ram_n18230, 
        p_wishbone_bd_ram_n18231, p_wishbone_bd_ram_n18232, 
        p_wishbone_bd_ram_n18233, p_wishbone_bd_ram_n18234, 
        p_wishbone_bd_ram_n18235, p_wishbone_bd_ram_n18236, 
        p_wishbone_bd_ram_n18237, p_wishbone_bd_ram_n18238, 
        p_wishbone_bd_ram_n18239, p_wishbone_bd_ram_n18240, 
        p_wishbone_bd_ram_n18241, p_wishbone_bd_ram_n18242, 
        p_wishbone_bd_ram_n18243, p_wishbone_bd_ram_n18244, 
        p_wishbone_bd_ram_n18245, p_wishbone_bd_ram_n18246, 
        p_wishbone_bd_ram_n18247, p_wishbone_bd_ram_n18248, 
        p_wishbone_bd_ram_n18249, p_wishbone_bd_ram_n18250, 
        p_wishbone_bd_ram_n18251, p_wishbone_bd_ram_n18252, 
        p_wishbone_bd_ram_n18253, p_wishbone_bd_ram_n18254, 
        p_wishbone_bd_ram_n18255, p_wishbone_bd_ram_n18256, 
        p_wishbone_bd_ram_n18257, p_wishbone_bd_ram_n18258, 
        p_wishbone_bd_ram_n18259, p_wishbone_bd_ram_n18260, 
        p_wishbone_bd_ram_n18261, p_wishbone_bd_ram_n18262, 
        p_wishbone_bd_ram_n18263, p_wishbone_bd_ram_n18264, 
        p_wishbone_bd_ram_n18265, p_wishbone_bd_ram_n18266, 
        p_wishbone_bd_ram_n18267, p_wishbone_bd_ram_n18268, 
        p_wishbone_bd_ram_n18269, p_wishbone_bd_ram_n18270, 
        p_wishbone_bd_ram_n18271, p_wishbone_bd_ram_n18272, 
        p_wishbone_bd_ram_n18273, p_wishbone_bd_ram_n18274, 
        p_wishbone_bd_ram_n18275, p_wishbone_bd_ram_n18276, 
        p_wishbone_bd_ram_n18277, p_wishbone_bd_ram_n18278, 
        p_wishbone_bd_ram_n18279, p_wishbone_bd_ram_n18280, 
        p_wishbone_bd_ram_n18281, p_wishbone_bd_ram_n18282, 
        p_wishbone_bd_ram_n18283, p_wishbone_bd_ram_n18284, 
        p_wishbone_bd_ram_n18285, p_wishbone_bd_ram_n18286, 
        p_wishbone_bd_ram_n18287, p_wishbone_bd_ram_n18288, 
        p_wishbone_bd_ram_n18289, p_wishbone_bd_ram_n18290, 
        p_wishbone_bd_ram_n18291, p_wishbone_bd_ram_n18292, 
        p_wishbone_bd_ram_n18293, p_wishbone_bd_ram_n18294, 
        p_wishbone_bd_ram_n18295, p_wishbone_bd_ram_n18296, 
        p_wishbone_bd_ram_n18297, p_wishbone_bd_ram_n18298, 
        p_wishbone_bd_ram_n18299, p_wishbone_bd_ram_n18300, 
        p_wishbone_bd_ram_n18301, p_wishbone_bd_ram_n18302, 
        p_wishbone_bd_ram_n18303, p_wishbone_bd_ram_n18304, 
        p_wishbone_bd_ram_n18305, p_wishbone_bd_ram_n18306, 
        p_wishbone_bd_ram_n18307, p_wishbone_bd_ram_n18308, 
        p_wishbone_bd_ram_n18309, p_wishbone_bd_ram_n18310, 
        p_wishbone_bd_ram_n18311, p_wishbone_bd_ram_n18312, 
        p_wishbone_bd_ram_n18313, p_wishbone_bd_ram_n18314, 
        p_wishbone_bd_ram_n18315, p_wishbone_bd_ram_n18316, 
        p_wishbone_bd_ram_n18317, p_wishbone_bd_ram_n18318, 
        p_wishbone_bd_ram_n18319, p_wishbone_bd_ram_n18320, 
        p_wishbone_bd_ram_n18321, p_wishbone_bd_ram_n18322, 
        p_wishbone_bd_ram_n18323, p_wishbone_bd_ram_n18324, 
        p_wishbone_bd_ram_n18325, p_wishbone_bd_ram_n18326, 
        p_wishbone_bd_ram_n18327, p_wishbone_bd_ram_n18328, 
        p_wishbone_bd_ram_n18329, p_wishbone_bd_ram_n18330, 
        p_wishbone_bd_ram_n18331, p_wishbone_bd_ram_n18332, 
        p_wishbone_bd_ram_n18333, p_wishbone_bd_ram_n18334, 
        p_wishbone_bd_ram_n18335, p_wishbone_bd_ram_n18336, 
        p_wishbone_bd_ram_n18337, p_wishbone_bd_ram_n18338, 
        p_wishbone_bd_ram_n18339, p_wishbone_bd_ram_n18340, 
        p_wishbone_bd_ram_n18341, p_wishbone_bd_ram_n18342, 
        p_wishbone_bd_ram_n18343, p_wishbone_bd_ram_n18344, 
        p_wishbone_bd_ram_n18345, p_wishbone_bd_ram_n18346, 
        p_wishbone_bd_ram_n18347, p_wishbone_bd_ram_n18348, 
        p_wishbone_bd_ram_n18349, p_wishbone_bd_ram_n18350, 
        p_wishbone_bd_ram_n18351, p_wishbone_bd_ram_n18352, 
        p_wishbone_bd_ram_n18353, p_wishbone_bd_ram_n18354, 
        p_wishbone_bd_ram_n18355, p_wishbone_bd_ram_n18356, 
        p_wishbone_bd_ram_n18357, p_wishbone_bd_ram_n18358, 
        p_wishbone_bd_ram_n18359, p_wishbone_bd_ram_n18360, 
        p_wishbone_bd_ram_n18361, p_wishbone_bd_ram_n18362, 
        p_wishbone_bd_ram_n18363, p_wishbone_bd_ram_n18364, 
        p_wishbone_bd_ram_n18365, p_wishbone_bd_ram_n18366, 
        p_wishbone_bd_ram_n18367, p_wishbone_bd_ram_n18368, 
        p_wishbone_bd_ram_n18369, p_wishbone_bd_ram_n18370, 
        p_wishbone_bd_ram_n18371, p_wishbone_bd_ram_n18372, 
        p_wishbone_bd_ram_n18373, p_wishbone_bd_ram_n18374, 
        p_wishbone_bd_ram_n18375, p_wishbone_bd_ram_n18376, 
        p_wishbone_bd_ram_n18377, p_wishbone_bd_ram_n18378, 
        p_wishbone_bd_ram_n18379, p_wishbone_bd_ram_n18380, 
        p_wishbone_bd_ram_n18381, p_wishbone_bd_ram_n18382, 
        p_wishbone_bd_ram_n18383, p_wishbone_bd_ram_n18384, 
        p_wishbone_bd_ram_n18385, p_wishbone_bd_ram_n18386, 
        p_wishbone_bd_ram_n18387, p_wishbone_bd_ram_n18388, 
        p_wishbone_bd_ram_n18389, p_wishbone_bd_ram_n18390, 
        p_wishbone_bd_ram_n18391, p_wishbone_bd_ram_n18392, 
        p_wishbone_bd_ram_n18393, p_wishbone_bd_ram_n18394, 
        p_wishbone_bd_ram_n18395, p_wishbone_bd_ram_n18396, 
        p_wishbone_bd_ram_n18397, p_wishbone_bd_ram_n18398, 
        p_wishbone_bd_ram_n18399, p_wishbone_bd_ram_n18400, 
        p_wishbone_bd_ram_n18401, p_wishbone_bd_ram_n18402, 
        p_wishbone_bd_ram_n18403, p_wishbone_bd_ram_n18404, 
        p_wishbone_bd_ram_n18405, p_wishbone_bd_ram_n18406, 
        p_wishbone_bd_ram_n18407, p_wishbone_bd_ram_n18408, 
        p_wishbone_bd_ram_n18409, p_wishbone_bd_ram_n18410, 
        p_wishbone_bd_ram_n18411, p_wishbone_bd_ram_n18412, 
        p_wishbone_bd_ram_n18413, p_wishbone_bd_ram_n18414, 
        p_wishbone_bd_ram_n18415, p_wishbone_bd_ram_n18416, 
        p_wishbone_bd_ram_n18417, p_wishbone_bd_ram_n18418, 
        p_wishbone_bd_ram_n18419, p_wishbone_bd_ram_n18420, 
        p_wishbone_bd_ram_n18421, p_wishbone_bd_ram_n18422, 
        p_wishbone_bd_ram_n18423, p_wishbone_bd_ram_n18424, 
        p_wishbone_bd_ram_n18425, p_wishbone_bd_ram_n18426, 
        p_wishbone_bd_ram_n18427, p_wishbone_bd_ram_n18428, 
        p_wishbone_bd_ram_n18429, p_wishbone_bd_ram_n18430, 
        p_wishbone_bd_ram_n18431, p_wishbone_bd_ram_n18432, 
        p_wishbone_bd_ram_n18433, p_wishbone_bd_ram_n18434, 
        p_wishbone_bd_ram_n18435, p_wishbone_bd_ram_n18436, 
        p_wishbone_bd_ram_n18437, p_wishbone_bd_ram_n18438, 
        p_wishbone_bd_ram_n18439, p_wishbone_bd_ram_n18440, 
        p_wishbone_bd_ram_n18441, p_wishbone_bd_ram_n18442, 
        p_wishbone_bd_ram_n18443, p_wishbone_bd_ram_n18444, 
        p_wishbone_bd_ram_n18445, p_wishbone_bd_ram_n18446, 
        p_wishbone_bd_ram_n18447, p_wishbone_bd_ram_n18448, 
        p_wishbone_bd_ram_n18449, p_wishbone_bd_ram_n18450, 
        p_wishbone_bd_ram_n18451, p_wishbone_bd_ram_n18452, 
        p_wishbone_bd_ram_n18453, p_wishbone_bd_ram_n18454, 
        p_wishbone_bd_ram_n18455, p_wishbone_bd_ram_n18456, 
        p_wishbone_bd_ram_n18457, p_wishbone_bd_ram_n18458, 
        p_wishbone_bd_ram_n18459, p_wishbone_bd_ram_n18460, 
        p_wishbone_bd_ram_n18461, p_wishbone_bd_ram_n18462, 
        p_wishbone_bd_ram_n18463, p_wishbone_bd_ram_n18464, 
        p_wishbone_bd_ram_n18465, p_wishbone_bd_ram_n18466, 
        p_wishbone_bd_ram_n18467, p_wishbone_bd_ram_n18468, 
        p_wishbone_bd_ram_n18469, p_wishbone_bd_ram_n18470, 
        p_wishbone_bd_ram_n18471, p_wishbone_bd_ram_n18472, 
        p_wishbone_bd_ram_n18473, p_wishbone_bd_ram_n18474, 
        p_wishbone_bd_ram_n18475, p_wishbone_bd_ram_n18476, 
        p_wishbone_bd_ram_n18477, p_wishbone_bd_ram_n18478, 
        p_wishbone_bd_ram_n18479, p_wishbone_bd_ram_n18480, 
        p_wishbone_bd_ram_n18481, p_wishbone_bd_ram_n18482, 
        p_wishbone_bd_ram_n18483, p_wishbone_bd_ram_n18484, 
        p_wishbone_bd_ram_n18485, p_wishbone_bd_ram_n18486, 
        p_wishbone_bd_ram_n18487, p_wishbone_bd_ram_n18488, 
        p_wishbone_bd_ram_n18489, p_wishbone_bd_ram_n18490, 
        p_wishbone_bd_ram_n18491, p_wishbone_bd_ram_n18492, 
        p_wishbone_bd_ram_n18493, p_wishbone_bd_ram_n18494, 
        p_wishbone_bd_ram_n18495, p_wishbone_bd_ram_n18496, 
        p_wishbone_bd_ram_n18497, p_wishbone_bd_ram_n18498, 
        p_wishbone_bd_ram_n18499, p_wishbone_bd_ram_n18500, 
        p_wishbone_bd_ram_n18501, p_wishbone_bd_ram_n18502, 
        p_wishbone_bd_ram_n18503, p_wishbone_bd_ram_n18504, 
        p_wishbone_bd_ram_n18505, p_wishbone_bd_ram_n18506, 
        p_wishbone_bd_ram_n18507, p_wishbone_bd_ram_n18508, 
        p_wishbone_bd_ram_n18509, p_wishbone_bd_ram_n18510, 
        p_wishbone_bd_ram_n18511, p_wishbone_bd_ram_n18512, 
        p_wishbone_bd_ram_n18513, p_wishbone_bd_ram_n18514, 
        p_wishbone_bd_ram_n18515, p_wishbone_bd_ram_n18516, 
        p_wishbone_bd_ram_n18517, p_wishbone_bd_ram_n18518, 
        p_wishbone_bd_ram_n18519, p_wishbone_bd_ram_n18520, 
        p_wishbone_bd_ram_n18521, p_wishbone_bd_ram_n18522, 
        p_wishbone_bd_ram_n18523, p_wishbone_bd_ram_n18524, 
        p_wishbone_bd_ram_n18525, p_wishbone_bd_ram_n18526, 
        p_wishbone_bd_ram_n18527, p_wishbone_bd_ram_n18528, 
        p_wishbone_bd_ram_n18529, p_wishbone_bd_ram_n18530, 
        p_wishbone_bd_ram_n18531, p_wishbone_bd_ram_n18532, 
        p_wishbone_bd_ram_n18533, p_wishbone_bd_ram_n18534, 
        p_wishbone_bd_ram_n18535, p_wishbone_bd_ram_n18536, 
        p_wishbone_bd_ram_n18537, p_wishbone_bd_ram_n18538, 
        p_wishbone_bd_ram_n18539, p_wishbone_bd_ram_n18540, 
        p_wishbone_bd_ram_n18541, p_wishbone_bd_ram_n18542, 
        p_wishbone_bd_ram_n18543, p_wishbone_bd_ram_n18544, 
        p_wishbone_bd_ram_n18545, p_wishbone_bd_ram_n18546, 
        p_wishbone_bd_ram_n18547, p_wishbone_bd_ram_n18548, 
        p_wishbone_bd_ram_n18549, p_wishbone_bd_ram_n18550, 
        p_wishbone_bd_ram_n18551, p_wishbone_bd_ram_n18552, 
        p_wishbone_bd_ram_n18553, p_wishbone_bd_ram_n18554, 
        p_wishbone_bd_ram_n18555, p_wishbone_bd_ram_n18556, 
        p_wishbone_bd_ram_n18557, p_wishbone_bd_ram_n18558, 
        p_wishbone_bd_ram_n18559, p_wishbone_bd_ram_n18560, 
        p_wishbone_bd_ram_n18561, p_wishbone_bd_ram_n18562, 
        p_wishbone_bd_ram_n18563, p_wishbone_bd_ram_n18564, 
        p_wishbone_bd_ram_n18565, p_wishbone_bd_ram_n18566, 
        p_wishbone_bd_ram_n18567, p_wishbone_bd_ram_n18568, 
        p_wishbone_bd_ram_n18569, p_wishbone_bd_ram_n18570, 
        p_wishbone_bd_ram_n18571, p_wishbone_bd_ram_n18572, 
        p_wishbone_bd_ram_n18573, p_wishbone_bd_ram_n18574, 
        p_wishbone_bd_ram_n18575, p_wishbone_bd_ram_n18576, 
        p_wishbone_bd_ram_n18577, p_wishbone_bd_ram_n18578, 
        p_wishbone_bd_ram_n18579, p_wishbone_bd_ram_n18580, 
        p_wishbone_bd_ram_n18581, p_wishbone_bd_ram_n18582, 
        p_wishbone_bd_ram_n18583, p_wishbone_bd_ram_n18584, 
        p_wishbone_bd_ram_n18585, p_wishbone_bd_ram_n18586, 
        p_wishbone_bd_ram_n18587, p_wishbone_bd_ram_n18588, 
        p_wishbone_bd_ram_n18589, p_wishbone_bd_ram_n18590, 
        p_wishbone_bd_ram_n18591, p_wishbone_bd_ram_n18592, 
        p_wishbone_bd_ram_n18593, p_wishbone_bd_ram_n18594, 
        p_wishbone_bd_ram_n18595, p_wishbone_bd_ram_n18596, 
        p_wishbone_bd_ram_n18597, p_wishbone_bd_ram_n18598, 
        p_wishbone_bd_ram_n18599, p_wishbone_bd_ram_n18600, 
        p_wishbone_bd_ram_n18601, p_wishbone_bd_ram_n18602, 
        p_wishbone_bd_ram_n18603, p_wishbone_bd_ram_n18604, 
        p_wishbone_bd_ram_n18605, p_wishbone_bd_ram_n18606, 
        p_wishbone_bd_ram_n18607, p_wishbone_bd_ram_n18608, 
        p_wishbone_bd_ram_n18609, p_wishbone_bd_ram_n18610, 
        p_wishbone_bd_ram_n18611, p_wishbone_bd_ram_n18612, 
        p_wishbone_bd_ram_n18613, p_wishbone_bd_ram_n18614, 
        p_wishbone_bd_ram_n18615, p_wishbone_bd_ram_n18616, 
        p_wishbone_bd_ram_n18617, p_wishbone_bd_ram_n18618, 
        p_wishbone_bd_ram_n18619, p_wishbone_bd_ram_n18620, 
        p_wishbone_bd_ram_n18621, p_wishbone_bd_ram_n18622, 
        p_wishbone_bd_ram_n18623, p_wishbone_bd_ram_n18624, 
        p_wishbone_bd_ram_n18625, p_wishbone_bd_ram_n18626, 
        p_wishbone_bd_ram_n18627, p_wishbone_bd_ram_n18628, 
        p_wishbone_bd_ram_n18629, p_wishbone_bd_ram_n18630, 
        p_wishbone_bd_ram_n18631, p_wishbone_bd_ram_n18632, 
        p_wishbone_bd_ram_n18633, p_wishbone_bd_ram_n18634, 
        p_wishbone_bd_ram_n18635, p_wishbone_bd_ram_n18636, 
        p_wishbone_bd_ram_n18637, p_wishbone_bd_ram_n18638, 
        p_wishbone_bd_ram_n18639, p_wishbone_bd_ram_n18640, 
        p_wishbone_bd_ram_n18641, p_wishbone_bd_ram_n18642, 
        p_wishbone_bd_ram_n18643, p_wishbone_bd_ram_n18644, 
        p_wishbone_bd_ram_n18645, p_wishbone_bd_ram_n18646, 
        p_wishbone_bd_ram_n18647, p_wishbone_bd_ram_n18648, 
        p_wishbone_bd_ram_n18649, p_wishbone_bd_ram_n18650, 
        p_wishbone_bd_ram_n18651, p_wishbone_bd_ram_n18652, 
        p_wishbone_bd_ram_n18653, p_wishbone_bd_ram_n18654, 
        p_wishbone_bd_ram_n18655, p_wishbone_bd_ram_n18656, 
        p_wishbone_bd_ram_n18657, p_wishbone_bd_ram_n18658, 
        p_wishbone_bd_ram_n18659, p_wishbone_bd_ram_n18660, 
        p_wishbone_bd_ram_n18661, p_wishbone_bd_ram_n18662, 
        p_wishbone_bd_ram_n18663, p_wishbone_bd_ram_n18664, 
        p_wishbone_bd_ram_n18665, p_wishbone_bd_ram_n18666, 
        p_wishbone_bd_ram_n18667, p_wishbone_bd_ram_n18668, 
        p_wishbone_bd_ram_n18669, p_wishbone_bd_ram_n18670, 
        p_wishbone_bd_ram_n18671, p_wishbone_bd_ram_n18672, 
        p_wishbone_bd_ram_n18673, p_wishbone_bd_ram_n18674, 
        p_wishbone_bd_ram_n18675, p_wishbone_bd_ram_n18676, 
        p_wishbone_bd_ram_n18677, p_wishbone_bd_ram_n18678, 
        p_wishbone_bd_ram_n18679, p_wishbone_bd_ram_n18680, 
        p_wishbone_bd_ram_n18681, p_wishbone_bd_ram_n18682, 
        p_wishbone_bd_ram_n18683, p_wishbone_bd_ram_n18684, 
        p_wishbone_bd_ram_n18685, p_wishbone_bd_ram_n18686, 
        p_wishbone_bd_ram_n18687, p_wishbone_bd_ram_n18688, 
        p_wishbone_bd_ram_n18689, p_wishbone_bd_ram_n18690, 
        p_wishbone_bd_ram_n18691, p_wishbone_bd_ram_n18692, 
        p_wishbone_bd_ram_n18693, p_wishbone_bd_ram_n18694, 
        p_wishbone_bd_ram_n18695, p_wishbone_bd_ram_n18696, 
        p_wishbone_bd_ram_n18697, p_wishbone_bd_ram_n18698, 
        p_wishbone_bd_ram_n18699, p_wishbone_bd_ram_n18700, 
        p_wishbone_bd_ram_n18701, p_wishbone_bd_ram_n18702, 
        p_wishbone_bd_ram_n18703, p_wishbone_bd_ram_n18704, 
        p_wishbone_bd_ram_n18705, p_wishbone_bd_ram_n18706, 
        p_wishbone_bd_ram_n18707, p_wishbone_bd_ram_n18708, 
        p_wishbone_bd_ram_n18709, p_wishbone_bd_ram_n18710, 
        p_wishbone_bd_ram_n18711, p_wishbone_bd_ram_n18712, 
        p_wishbone_bd_ram_n18713, p_wishbone_bd_ram_n18714, 
        p_wishbone_bd_ram_n18715, p_wishbone_bd_ram_n18716, 
        p_wishbone_bd_ram_n18717, p_wishbone_bd_ram_n18718, 
        p_wishbone_bd_ram_n18719, p_wishbone_bd_ram_n18720, 
        p_wishbone_bd_ram_n18721, p_wishbone_bd_ram_n18722, 
        p_wishbone_bd_ram_n18723, p_wishbone_bd_ram_n18724, 
        p_wishbone_bd_ram_n18725, p_wishbone_bd_ram_n18726, 
        p_wishbone_bd_ram_n18727, p_wishbone_bd_ram_n18728, 
        p_wishbone_bd_ram_n18729, p_wishbone_bd_ram_n18730, 
        p_wishbone_bd_ram_n18731, p_wishbone_bd_ram_n18732, 
        p_wishbone_bd_ram_n18733, p_wishbone_bd_ram_n18734, 
        p_wishbone_bd_ram_n18735, p_wishbone_bd_ram_n18736, 
        p_wishbone_bd_ram_n18737, p_wishbone_bd_ram_n18738, 
        p_wishbone_bd_ram_n18739, p_wishbone_bd_ram_n18740, 
        p_wishbone_bd_ram_n18741, p_wishbone_bd_ram_n18742, 
        p_wishbone_bd_ram_n18743, p_wishbone_bd_ram_n18744, 
        p_wishbone_bd_ram_n18745, p_wishbone_bd_ram_n18746, 
        p_wishbone_bd_ram_n18747, p_wishbone_bd_ram_n18748, 
        p_wishbone_bd_ram_n18749, p_wishbone_bd_ram_n18750, 
        p_wishbone_bd_ram_n18751, p_wishbone_bd_ram_n18752, 
        p_wishbone_bd_ram_n18753, p_wishbone_bd_ram_n18754, 
        p_wishbone_bd_ram_n18755, p_wishbone_bd_ram_n18756, 
        p_wishbone_bd_ram_n18757, p_wishbone_bd_ram_n18758, 
        p_wishbone_bd_ram_n18759, p_wishbone_bd_ram_n18760, 
        p_wishbone_bd_ram_n18761, p_wishbone_bd_ram_n18762, 
        p_wishbone_bd_ram_n18763, p_wishbone_bd_ram_n18764, 
        p_wishbone_bd_ram_n18765, p_wishbone_bd_ram_n18766, 
        p_wishbone_bd_ram_n18767, p_wishbone_bd_ram_n18768, 
        p_wishbone_bd_ram_n18769, p_wishbone_bd_ram_n18770, 
        p_wishbone_bd_ram_n18771, p_wishbone_bd_ram_n18772, 
        p_wishbone_bd_ram_n18773, p_wishbone_bd_ram_n18774, 
        p_wishbone_bd_ram_n18775, p_wishbone_bd_ram_n18776, 
        p_wishbone_bd_ram_n18777, p_wishbone_bd_ram_n18778, 
        p_wishbone_bd_ram_n18779, p_wishbone_bd_ram_n18780, 
        p_wishbone_bd_ram_n18781, p_wishbone_bd_ram_n18782, 
        p_wishbone_bd_ram_n18783, p_wishbone_bd_ram_n18784, 
        p_wishbone_bd_ram_n18785, p_wishbone_bd_ram_n18786, 
        p_wishbone_bd_ram_n18787, p_wishbone_bd_ram_n18788, 
        p_wishbone_bd_ram_n18789, p_wishbone_bd_ram_n18790, 
        p_wishbone_bd_ram_n18791, p_wishbone_bd_ram_n18792, 
        p_wishbone_bd_ram_n18793, p_wishbone_bd_ram_n18794, 
        p_wishbone_bd_ram_n18795, p_wishbone_bd_ram_n18796, 
        p_wishbone_bd_ram_n18797, p_wishbone_bd_ram_n18798, 
        p_wishbone_bd_ram_n18799, p_wishbone_bd_ram_n18800, 
        p_wishbone_bd_ram_n18801, p_wishbone_bd_ram_n18802, 
        p_wishbone_bd_ram_n18803, p_wishbone_bd_ram_n18804, 
        p_wishbone_bd_ram_n18805, p_wishbone_bd_ram_n18806, 
        p_wishbone_bd_ram_n18807, p_wishbone_bd_ram_n18808, 
        p_wishbone_bd_ram_n18809, p_wishbone_bd_ram_n18810, 
        p_wishbone_bd_ram_n18811, p_wishbone_bd_ram_n18812, 
        p_wishbone_bd_ram_n18813, p_wishbone_bd_ram_n18814, 
        p_wishbone_bd_ram_n18815, p_wishbone_bd_ram_n18816, 
        p_wishbone_bd_ram_n18817, p_wishbone_bd_ram_n18818, 
        p_wishbone_bd_ram_n18819, p_wishbone_bd_ram_n18820, 
        p_wishbone_bd_ram_n18821, p_wishbone_bd_ram_n18822, 
        p_wishbone_bd_ram_n18823, p_wishbone_bd_ram_n18824, 
        p_wishbone_bd_ram_n18825, p_wishbone_bd_ram_n18826, 
        p_wishbone_bd_ram_n18827, p_wishbone_bd_ram_n18828, 
        p_wishbone_bd_ram_n18829, p_wishbone_bd_ram_n18830, 
        p_wishbone_bd_ram_n18831, p_wishbone_bd_ram_n18832, 
        p_wishbone_bd_ram_n18833, p_wishbone_bd_ram_n18834, 
        p_wishbone_bd_ram_n18835, p_wishbone_bd_ram_n18836, 
        p_wishbone_bd_ram_n18837, p_wishbone_bd_ram_n18838, 
        p_wishbone_bd_ram_n18839, p_wishbone_bd_ram_n18840, 
        p_wishbone_bd_ram_n18841, p_wishbone_bd_ram_n18842, 
        p_wishbone_bd_ram_n18843, p_wishbone_bd_ram_n18844, 
        p_wishbone_bd_ram_n18845, p_wishbone_bd_ram_n18846, 
        p_wishbone_bd_ram_n18847, p_wishbone_bd_ram_n18848, 
        p_wishbone_bd_ram_n18849, p_wishbone_bd_ram_n18850, 
        p_wishbone_bd_ram_n18851, p_wishbone_bd_ram_n18852, 
        p_wishbone_bd_ram_n18853, p_wishbone_bd_ram_n18854, 
        p_wishbone_bd_ram_n18855, p_wishbone_bd_ram_n18856, 
        p_wishbone_bd_ram_n18857, p_wishbone_bd_ram_n18858, 
        p_wishbone_bd_ram_n18859, p_wishbone_bd_ram_n18860, 
        p_wishbone_bd_ram_n18861, p_wishbone_bd_ram_n18862, 
        p_wishbone_bd_ram_n18863, p_wishbone_bd_ram_n18864, 
        p_wishbone_bd_ram_n18865, p_wishbone_bd_ram_n18866, 
        p_wishbone_bd_ram_n18867, p_wishbone_bd_ram_n18868, 
        p_wishbone_bd_ram_n18869, p_wishbone_bd_ram_n18870, 
        p_wishbone_bd_ram_n18871, p_wishbone_bd_ram_n18872, 
        p_wishbone_bd_ram_n18873, p_wishbone_bd_ram_n18874, 
        p_wishbone_bd_ram_n18875, p_wishbone_bd_ram_n18876, 
        p_wishbone_bd_ram_n18877, p_wishbone_bd_ram_n18878, 
        p_wishbone_bd_ram_n18879, p_wishbone_bd_ram_n18880, 
        p_wishbone_bd_ram_n18881, p_wishbone_bd_ram_n18882, 
        p_wishbone_bd_ram_n18883, p_wishbone_bd_ram_n18884, 
        p_wishbone_bd_ram_n18885, p_wishbone_bd_ram_n18886, 
        p_wishbone_bd_ram_n18887, p_wishbone_bd_ram_n18888, 
        p_wishbone_bd_ram_n18889, p_wishbone_bd_ram_n18890, 
        p_wishbone_bd_ram_n18891, p_wishbone_bd_ram_n18892, 
        p_wishbone_bd_ram_n18893, p_wishbone_bd_ram_n18894, 
        p_wishbone_bd_ram_n18895, p_wishbone_bd_ram_n18896, 
        p_wishbone_bd_ram_n18897, p_wishbone_bd_ram_n18898, 
        p_wishbone_bd_ram_n18899, p_wishbone_bd_ram_n18900, 
        p_wishbone_bd_ram_n18901, p_wishbone_bd_ram_n18902, 
        p_wishbone_bd_ram_n18903, p_wishbone_bd_ram_n18904, 
        p_wishbone_bd_ram_n18905, p_wishbone_bd_ram_n18906, 
        p_wishbone_bd_ram_n18907, p_wishbone_bd_ram_n18908, 
        p_wishbone_bd_ram_n18909, p_wishbone_bd_ram_n18910, 
        p_wishbone_bd_ram_n18911, p_wishbone_bd_ram_n18912, 
        p_wishbone_bd_ram_n18913, p_wishbone_bd_ram_n18914, 
        p_wishbone_bd_ram_n18915, p_wishbone_bd_ram_n18916, 
        p_wishbone_bd_ram_n18917, p_wishbone_bd_ram_n18918, 
        p_wishbone_bd_ram_n18919, p_wishbone_bd_ram_n18920, 
        p_wishbone_bd_ram_n18921, p_wishbone_bd_ram_n18922, 
        p_wishbone_bd_ram_n18923, p_wishbone_bd_ram_n18924, 
        p_wishbone_bd_ram_n18925, p_wishbone_bd_ram_n18926, 
        p_wishbone_bd_ram_n18927, p_wishbone_bd_ram_n18928, 
        p_wishbone_bd_ram_n18929, p_wishbone_bd_ram_n18930, 
        p_wishbone_bd_ram_n18931, p_wishbone_bd_ram_n18932, 
        p_wishbone_bd_ram_n18933, p_wishbone_bd_ram_n18934, 
        p_wishbone_bd_ram_n18935, p_wishbone_bd_ram_n18936, 
        p_wishbone_bd_ram_n18937, p_wishbone_bd_ram_n18938, 
        p_wishbone_bd_ram_n18939, p_wishbone_bd_ram_n18940, 
        p_wishbone_bd_ram_n18941, p_wishbone_bd_ram_n18942, 
        p_wishbone_bd_ram_n18943, p_wishbone_bd_ram_n18944, 
        p_wishbone_bd_ram_n18945, p_wishbone_bd_ram_n18946, 
        p_wishbone_bd_ram_n18947, p_wishbone_bd_ram_n18948, 
        p_wishbone_bd_ram_n18949, p_wishbone_bd_ram_n18950, 
        p_wishbone_bd_ram_n18951, p_wishbone_bd_ram_n18952, 
        p_wishbone_bd_ram_n18953, p_wishbone_bd_ram_n18954, 
        p_wishbone_bd_ram_n18955, p_wishbone_bd_ram_n18956, 
        p_wishbone_bd_ram_n18957, p_wishbone_bd_ram_n18958, 
        p_wishbone_bd_ram_n18959, p_wishbone_bd_ram_n18960, 
        p_wishbone_bd_ram_n18961, p_wishbone_bd_ram_n18962, 
        p_wishbone_bd_ram_n18963, p_wishbone_bd_ram_n18964, 
        p_wishbone_bd_ram_n18965, p_wishbone_bd_ram_n18966, 
        p_wishbone_bd_ram_n18967, p_wishbone_bd_ram_n18968, 
        p_wishbone_bd_ram_n18969, p_wishbone_bd_ram_n18970, 
        p_wishbone_bd_ram_n18971, p_wishbone_bd_ram_n18972, 
        p_wishbone_bd_ram_n18973, p_wishbone_bd_ram_n18974, 
        p_wishbone_bd_ram_n18975, p_wishbone_bd_ram_n18976, 
        p_wishbone_bd_ram_n18977, p_wishbone_bd_ram_n18978, 
        p_wishbone_bd_ram_n18979, p_wishbone_bd_ram_n18980, 
        p_wishbone_bd_ram_n18981, p_wishbone_bd_ram_n18982, 
        p_wishbone_bd_ram_n18983, p_wishbone_bd_ram_n18984, 
        p_wishbone_bd_ram_n18985, p_wishbone_bd_ram_n18986, 
        p_wishbone_bd_ram_n18987, p_wishbone_bd_ram_n18988, 
        p_wishbone_bd_ram_n18989, p_wishbone_bd_ram_n18990, 
        p_wishbone_bd_ram_n18991, p_wishbone_bd_ram_n18992, 
        p_wishbone_bd_ram_n18993, p_wishbone_bd_ram_n18994, 
        p_wishbone_bd_ram_n18995, p_wishbone_bd_ram_n18996, 
        p_wishbone_bd_ram_n18997, p_wishbone_bd_ram_n18998, 
        p_wishbone_bd_ram_n18999, p_wishbone_bd_ram_n19000, 
        p_wishbone_bd_ram_n19001, p_wishbone_bd_ram_n19002, 
        p_wishbone_bd_ram_n19003, p_wishbone_bd_ram_n19004, 
        p_wishbone_bd_ram_n19005, p_wishbone_bd_ram_n19006, 
        p_wishbone_bd_ram_n19007, p_wishbone_bd_ram_n19008, 
        p_wishbone_bd_ram_n19009, p_wishbone_bd_ram_n19010, 
        p_wishbone_bd_ram_n19011, p_wishbone_bd_ram_n19012, 
        p_wishbone_bd_ram_n19013, p_wishbone_bd_ram_n19014, 
        p_wishbone_bd_ram_n19015, p_wishbone_bd_ram_n19016, 
        p_wishbone_bd_ram_n19017, p_wishbone_bd_ram_n19018, 
        p_wishbone_bd_ram_n19019, p_wishbone_bd_ram_n19020, 
        p_wishbone_bd_ram_n19021, p_wishbone_bd_ram_n19022, 
        p_wishbone_bd_ram_n19023, p_wishbone_bd_ram_n19024, 
        p_wishbone_bd_ram_n19025, p_wishbone_bd_ram_n19026, 
        p_wishbone_bd_ram_n19027, p_wishbone_bd_ram_n19028, 
        p_wishbone_bd_ram_n19029, p_wishbone_bd_ram_n19030, 
        p_wishbone_bd_ram_n19031, p_wishbone_bd_ram_n19032, 
        p_wishbone_bd_ram_n19033, p_wishbone_bd_ram_n19034, 
        p_wishbone_bd_ram_n19035, p_wishbone_bd_ram_n19036, 
        p_wishbone_bd_ram_n19037, p_wishbone_bd_ram_n19038, 
        p_wishbone_bd_ram_n19039, p_wishbone_bd_ram_n19040, 
        p_wishbone_bd_ram_n19041, p_wishbone_bd_ram_n19042, 
        p_wishbone_bd_ram_n19043, p_wishbone_bd_ram_n19044, 
        p_wishbone_bd_ram_n19045, p_wishbone_bd_ram_n19046, 
        p_wishbone_bd_ram_n19047, p_wishbone_bd_ram_n19048, 
        p_wishbone_bd_ram_n19049, p_wishbone_bd_ram_n19050, 
        p_wishbone_bd_ram_n19051, p_wishbone_bd_ram_n19052, 
        p_wishbone_bd_ram_n19053, p_wishbone_bd_ram_n19054, 
        p_wishbone_bd_ram_n19055, p_wishbone_bd_ram_n19056, 
        p_wishbone_bd_ram_n19057, p_wishbone_bd_ram_n19058, 
        p_wishbone_bd_ram_n19059, p_wishbone_bd_ram_n19060, 
        p_wishbone_bd_ram_n19061, p_wishbone_bd_ram_n19062, 
        p_wishbone_bd_ram_n19063, p_wishbone_bd_ram_n19064, 
        p_wishbone_bd_ram_n19065, p_wishbone_bd_ram_n19066, 
        p_wishbone_bd_ram_n19067, p_wishbone_bd_ram_n19068, 
        p_wishbone_bd_ram_n19069, p_wishbone_bd_ram_n19070, 
        p_wishbone_bd_ram_n19071, p_wishbone_bd_ram_n19072, 
        p_wishbone_bd_ram_n19073, p_wishbone_bd_ram_n19074, 
        p_wishbone_bd_ram_n19075, p_wishbone_bd_ram_n19076, 
        p_wishbone_bd_ram_n19077, p_wishbone_bd_ram_n19078, 
        p_wishbone_bd_ram_n19079, p_wishbone_bd_ram_n19080, 
        p_wishbone_bd_ram_n19081, p_wishbone_bd_ram_n19082, 
        p_wishbone_bd_ram_n19083, p_wishbone_bd_ram_n19084, 
        p_wishbone_bd_ram_n19085, p_wishbone_bd_ram_n19086, 
        p_wishbone_bd_ram_n19087, p_wishbone_bd_ram_n19088, 
        p_wishbone_bd_ram_n19089, p_wishbone_bd_ram_n19090, 
        p_wishbone_bd_ram_n19091, p_wishbone_bd_ram_n19092, 
        p_wishbone_bd_ram_n19093, p_wishbone_bd_ram_n19094, 
        p_wishbone_bd_ram_n19095, p_wishbone_bd_ram_n19096, 
        p_wishbone_bd_ram_n19097, p_wishbone_bd_ram_n19098, 
        p_wishbone_bd_ram_n19099, p_wishbone_bd_ram_n19100, 
        p_wishbone_bd_ram_n19101, p_wishbone_bd_ram_n19102, 
        p_wishbone_bd_ram_n19103, p_wishbone_bd_ram_n19104, 
        p_wishbone_bd_ram_n19105, p_wishbone_bd_ram_n19106, 
        p_wishbone_bd_ram_n19107, p_wishbone_bd_ram_n19108, 
        p_wishbone_bd_ram_n19109, p_wishbone_bd_ram_n19110, 
        p_wishbone_bd_ram_n19111, p_wishbone_bd_ram_n19112, 
        p_wishbone_bd_ram_n19113, p_wishbone_bd_ram_n19114, 
        p_wishbone_bd_ram_n19115, p_wishbone_bd_ram_n19116, 
        p_wishbone_bd_ram_n19117, p_wishbone_bd_ram_n19118, 
        p_wishbone_bd_ram_n19119, p_wishbone_bd_ram_n19120, 
        p_wishbone_bd_ram_n19121, p_wishbone_bd_ram_n19122, 
        p_wishbone_bd_ram_n19123, p_wishbone_bd_ram_n19124, 
        p_wishbone_bd_ram_n19125, p_wishbone_bd_ram_n19126, 
        p_wishbone_bd_ram_n19127, p_wishbone_bd_ram_n19128, 
        p_wishbone_bd_ram_n19129, p_wishbone_bd_ram_n19130, 
        p_wishbone_bd_ram_n19131, p_wishbone_bd_ram_n19132, 
        p_wishbone_bd_ram_n19133, p_wishbone_bd_ram_n19134, 
        p_wishbone_bd_ram_n19135, p_wishbone_bd_ram_n19136, 
        p_wishbone_bd_ram_n19137, p_wishbone_bd_ram_n19138, 
        p_wishbone_bd_ram_n19139, p_wishbone_bd_ram_n19140, 
        p_wishbone_bd_ram_n19141, p_wishbone_bd_ram_n19142, 
        p_wishbone_bd_ram_n19143, p_wishbone_bd_ram_n19144, 
        p_wishbone_bd_ram_n19145, p_wishbone_bd_ram_n19146, 
        p_wishbone_bd_ram_n19147, p_wishbone_bd_ram_n19148, 
        p_wishbone_bd_ram_n19149, p_wishbone_bd_ram_n19150, 
        p_wishbone_bd_ram_n19151, p_wishbone_bd_ram_n19152, 
        p_wishbone_bd_ram_n19153, p_wishbone_bd_ram_n19154, 
        p_wishbone_bd_ram_n19155, p_wishbone_bd_ram_n19156, 
        p_wishbone_bd_ram_n19157, p_wishbone_bd_ram_n19158, 
        p_wishbone_bd_ram_n19159, p_wishbone_bd_ram_n19160, 
        p_wishbone_bd_ram_n19161, p_wishbone_bd_ram_n19162, 
        p_wishbone_bd_ram_n19163, p_wishbone_bd_ram_n19164, 
        p_wishbone_bd_ram_n19165, p_wishbone_bd_ram_n19166, 
        p_wishbone_bd_ram_n19167, p_wishbone_bd_ram_n19168, 
        p_wishbone_bd_ram_n19169, p_wishbone_bd_ram_n19170, 
        p_wishbone_bd_ram_n19171, p_wishbone_bd_ram_n19172, 
        p_wishbone_bd_ram_n19173, p_wishbone_bd_ram_n19174, 
        p_wishbone_bd_ram_n19175, p_wishbone_bd_ram_n19176, 
        p_wishbone_bd_ram_n19177, p_wishbone_bd_ram_n19178, 
        p_wishbone_bd_ram_n19179, p_wishbone_bd_ram_n19180, 
        p_wishbone_bd_ram_n19181, p_wishbone_bd_ram_n19182, 
        p_wishbone_bd_ram_n19183, p_wishbone_bd_ram_n19184, 
        p_wishbone_bd_ram_n19185, p_wishbone_bd_ram_n19186, 
        p_wishbone_bd_ram_n19187, p_wishbone_bd_ram_n19188, 
        p_wishbone_bd_ram_n19189, p_wishbone_bd_ram_n19190, 
        p_wishbone_bd_ram_n19191, p_wishbone_bd_ram_n19192, 
        p_wishbone_bd_ram_n19193, p_wishbone_bd_ram_n19194, 
        p_wishbone_bd_ram_n19195, p_wishbone_bd_ram_n19196, 
        p_wishbone_bd_ram_n19197, p_wishbone_bd_ram_n19198, 
        p_wishbone_bd_ram_n19199, p_wishbone_bd_ram_n19200, 
        p_wishbone_bd_ram_n19201, p_wishbone_bd_ram_n19202, 
        p_wishbone_bd_ram_n19203, p_wishbone_bd_ram_n19204, 
        p_wishbone_bd_ram_n19205, p_wishbone_bd_ram_n19206, 
        p_wishbone_bd_ram_n19207, p_wishbone_bd_ram_n19208, 
        p_wishbone_bd_ram_n19209, p_wishbone_bd_ram_n19210, 
        p_wishbone_bd_ram_n19211, p_wishbone_bd_ram_n19212, 
        p_wishbone_bd_ram_n19213, p_wishbone_bd_ram_n19214, 
        p_wishbone_bd_ram_n19215, p_wishbone_bd_ram_n19216, 
        p_wishbone_bd_ram_n19217, p_wishbone_bd_ram_n19218, 
        p_wishbone_bd_ram_n19219, p_wishbone_bd_ram_n19220, 
        p_wishbone_bd_ram_n19221, p_wishbone_bd_ram_n19222, 
        p_wishbone_bd_ram_n19223, p_wishbone_bd_ram_n19224, 
        p_wishbone_bd_ram_n19225, p_wishbone_bd_ram_n19226, 
        p_wishbone_bd_ram_n19227, p_wishbone_bd_ram_n19228, 
        p_wishbone_bd_ram_n19229, p_wishbone_bd_ram_n19230, 
        p_wishbone_bd_ram_n19231, p_wishbone_bd_ram_n19232, 
        p_wishbone_bd_ram_n19233, p_wishbone_bd_ram_n19234, 
        p_wishbone_bd_ram_n19235, p_wishbone_bd_ram_n19236, 
        p_wishbone_bd_ram_n19237, p_wishbone_bd_ram_n19238, 
        p_wishbone_bd_ram_n19239, p_wishbone_bd_ram_n19240, 
        p_wishbone_bd_ram_n19241, p_wishbone_bd_ram_n19242, 
        p_wishbone_bd_ram_n19243, p_wishbone_bd_ram_n19244, 
        p_wishbone_bd_ram_n19245, p_wishbone_bd_ram_n19246, 
        p_wishbone_bd_ram_n19247, p_wishbone_bd_ram_n19248, 
        p_wishbone_bd_ram_n19249, p_wishbone_bd_ram_n19250, 
        p_wishbone_bd_ram_n19251, p_wishbone_bd_ram_n19252, 
        p_wishbone_bd_ram_n19253, p_wishbone_bd_ram_n19254, 
        p_wishbone_bd_ram_n19255, p_wishbone_bd_ram_n19256, 
        p_wishbone_bd_ram_n19257, p_wishbone_bd_ram_n19258, 
        p_wishbone_bd_ram_n19259, p_wishbone_bd_ram_n19260, 
        p_wishbone_bd_ram_n19261, p_wishbone_bd_ram_n19262, 
        p_wishbone_bd_ram_n19263, p_wishbone_bd_ram_n19264, 
        p_wishbone_bd_ram_n19265, p_wishbone_bd_ram_n19266, 
        p_wishbone_bd_ram_n19267, p_wishbone_bd_ram_n19268, 
        p_wishbone_bd_ram_n19269, p_wishbone_bd_ram_n19270, 
        p_wishbone_bd_ram_n19271, p_wishbone_bd_ram_n19272, 
        p_wishbone_bd_ram_n19273, p_wishbone_bd_ram_n19274, 
        p_wishbone_bd_ram_n19275, p_wishbone_bd_ram_n19276, 
        p_wishbone_bd_ram_n19277, p_wishbone_bd_ram_n19278, 
        p_wishbone_bd_ram_n19279, p_wishbone_bd_ram_n19280, 
        p_wishbone_bd_ram_n19281, p_wishbone_bd_ram_n19282, 
        p_wishbone_bd_ram_n19283, p_wishbone_bd_ram_n19284, 
        p_wishbone_bd_ram_n19285, p_wishbone_bd_ram_n19286, 
        p_wishbone_bd_ram_n19287, p_wishbone_bd_ram_n19288, 
        p_wishbone_bd_ram_n19289, p_wishbone_bd_ram_n19290, 
        p_wishbone_bd_ram_n19291, p_wishbone_bd_ram_n19292, 
        p_wishbone_bd_ram_n19293, p_wishbone_bd_ram_n19294, 
        p_wishbone_bd_ram_n19295, p_wishbone_bd_ram_n19296, 
        p_wishbone_bd_ram_n19297, p_wishbone_bd_ram_n19298, 
        p_wishbone_bd_ram_n19299, p_wishbone_bd_ram_n19300, 
        p_wishbone_bd_ram_n19301, p_wishbone_bd_ram_n19302, 
        p_wishbone_bd_ram_n19303, p_wishbone_bd_ram_n19304, 
        p_wishbone_bd_ram_n19305, p_wishbone_bd_ram_n19306, 
        p_wishbone_bd_ram_n19307, p_wishbone_bd_ram_n19308, 
        p_wishbone_bd_ram_n19309, p_wishbone_bd_ram_n19310, 
        p_wishbone_bd_ram_n19311, p_wishbone_bd_ram_n19312, 
        p_wishbone_bd_ram_n19313, p_wishbone_bd_ram_n19314, 
        p_wishbone_bd_ram_n19315, p_wishbone_bd_ram_n19316, 
        p_wishbone_bd_ram_n19317, p_wishbone_bd_ram_n19318, 
        p_wishbone_bd_ram_n19319, p_wishbone_bd_ram_n19320, 
        p_wishbone_bd_ram_n19321, p_wishbone_bd_ram_n19322, 
        p_wishbone_bd_ram_n19323, p_wishbone_bd_ram_n19324, 
        p_wishbone_bd_ram_n19325, p_wishbone_bd_ram_n19326, 
        p_wishbone_bd_ram_n19327, p_wishbone_bd_ram_n19328, 
        p_wishbone_bd_ram_n19329, p_wishbone_bd_ram_n19330, 
        p_wishbone_bd_ram_n19331, p_wishbone_bd_ram_n19332, 
        p_wishbone_bd_ram_n19333, p_wishbone_bd_ram_n19334, 
        p_wishbone_bd_ram_n19335, p_wishbone_bd_ram_n19336, 
        p_wishbone_bd_ram_n19337, p_wishbone_bd_ram_n19338, 
        p_wishbone_bd_ram_n19339, p_wishbone_bd_ram_n19340, 
        p_wishbone_bd_ram_n19341, p_wishbone_bd_ram_n19342, 
        p_wishbone_bd_ram_n19343, p_wishbone_bd_ram_n19344, 
        p_wishbone_bd_ram_n19345, p_wishbone_bd_ram_n19346, 
        p_wishbone_bd_ram_n19347, p_wishbone_bd_ram_n19348, 
        p_wishbone_bd_ram_n19349, p_wishbone_bd_ram_n19350, 
        p_wishbone_bd_ram_n19351, p_wishbone_bd_ram_n19352, 
        p_wishbone_bd_ram_n19353, p_wishbone_bd_ram_n19354, 
        p_wishbone_bd_ram_n19355, p_wishbone_bd_ram_n19356, 
        p_wishbone_bd_ram_n19357, p_wishbone_bd_ram_n19358, 
        p_wishbone_bd_ram_n19359, p_wishbone_bd_ram_n19360, 
        p_wishbone_bd_ram_n19361, p_wishbone_bd_ram_n19362, 
        p_wishbone_bd_ram_n19363, p_wishbone_bd_ram_n19364, 
        p_wishbone_bd_ram_n19365, p_wishbone_bd_ram_n19366, 
        p_wishbone_bd_ram_n19367, p_wishbone_bd_ram_n19368, 
        p_wishbone_bd_ram_n19369, p_wishbone_bd_ram_n19370, 
        p_wishbone_bd_ram_n19371, p_wishbone_bd_ram_n19372, 
        p_wishbone_bd_ram_n19373, p_wishbone_bd_ram_n19374, 
        p_wishbone_bd_ram_n19375, p_wishbone_bd_ram_n19376, 
        p_wishbone_bd_ram_n19377, p_wishbone_bd_ram_n19378, 
        p_wishbone_bd_ram_n19379, p_wishbone_bd_ram_n19380, 
        p_wishbone_bd_ram_n19381, p_wishbone_bd_ram_n19382, 
        p_wishbone_bd_ram_n19383, p_wishbone_bd_ram_n19384, 
        p_wishbone_bd_ram_n19385, p_wishbone_bd_ram_n19386, 
        p_wishbone_bd_ram_n19387, p_wishbone_bd_ram_n19388, 
        p_wishbone_bd_ram_n19389, p_wishbone_bd_ram_n19390, 
        p_wishbone_bd_ram_n19391, p_wishbone_bd_ram_n19392, 
        p_wishbone_bd_ram_n19393, p_wishbone_bd_ram_n19394, 
        p_wishbone_bd_ram_n19395, p_wishbone_bd_ram_n19396, 
        p_wishbone_bd_ram_n19397, p_wishbone_bd_ram_n19398, 
        p_wishbone_bd_ram_n19399, p_wishbone_bd_ram_n19400, 
        p_wishbone_bd_ram_n19401, p_wishbone_bd_ram_n19402, 
        p_wishbone_bd_ram_n19403, p_wishbone_bd_ram_n19404, 
        p_wishbone_bd_ram_n19405, p_wishbone_bd_ram_n19406, 
        p_wishbone_bd_ram_n19407, p_wishbone_bd_ram_n19408, 
        p_wishbone_bd_ram_n19409, p_wishbone_bd_ram_n19410, 
        p_wishbone_bd_ram_n19411, p_wishbone_bd_ram_n19412, 
        p_wishbone_bd_ram_n19413, p_wishbone_bd_ram_n19414, 
        p_wishbone_bd_ram_n19415, p_wishbone_bd_ram_n19416, 
        p_wishbone_bd_ram_n19417, p_wishbone_bd_ram_n19418, 
        p_wishbone_bd_ram_n19419, p_wishbone_bd_ram_n19420, 
        p_wishbone_bd_ram_n19421, p_wishbone_bd_ram_n19422, 
        p_wishbone_bd_ram_n19423, p_wishbone_bd_ram_n19424, 
        p_wishbone_bd_ram_n19425, p_wishbone_bd_ram_n19426, 
        p_wishbone_bd_ram_n19427, p_wishbone_bd_ram_n19428, 
        p_wishbone_bd_ram_n19429, p_wishbone_bd_ram_n19430, 
        p_wishbone_bd_ram_n19431, p_wishbone_bd_ram_n19432, 
        p_wishbone_bd_ram_n19433, p_wishbone_bd_ram_n19434, 
        p_wishbone_bd_ram_n19435, p_wishbone_bd_ram_n19436, 
        p_wishbone_bd_ram_n19437, p_wishbone_bd_ram_n19438, 
        p_wishbone_bd_ram_n19439, p_wishbone_bd_ram_n19440, 
        p_wishbone_bd_ram_n19441, p_wishbone_bd_ram_n19442, 
        p_wishbone_bd_ram_n19443, p_wishbone_bd_ram_n19444, 
        p_wishbone_bd_ram_n19445, p_wishbone_bd_ram_n19446, 
        p_wishbone_bd_ram_n19447, p_wishbone_bd_ram_n19448, 
        p_wishbone_bd_ram_n19449, p_wishbone_bd_ram_n19450, 
        p_wishbone_bd_ram_n19451, p_wishbone_bd_ram_n19452, 
        p_wishbone_bd_ram_n19453, p_wishbone_bd_ram_n19454, 
        p_wishbone_bd_ram_n19455, p_wishbone_bd_ram_n19456, 
        p_wishbone_bd_ram_n19457, p_wishbone_bd_ram_n19458, 
        p_wishbone_bd_ram_n19459, p_wishbone_bd_ram_n19460, 
        p_wishbone_bd_ram_n19461, p_wishbone_bd_ram_n19462, 
        p_wishbone_bd_ram_n19463, p_wishbone_bd_ram_n19464, 
        p_wishbone_bd_ram_n19465, p_wishbone_bd_ram_n19466, 
        p_wishbone_bd_ram_n19467, p_wishbone_bd_ram_n19468, 
        p_wishbone_bd_ram_n19469, p_wishbone_bd_ram_n19470, 
        p_wishbone_bd_ram_n19471, p_wishbone_bd_ram_n19472, 
        p_wishbone_bd_ram_n19473, p_wishbone_bd_ram_n19474, 
        p_wishbone_bd_ram_n19475, p_wishbone_bd_ram_n19476, 
        p_wishbone_bd_ram_n19477, p_wishbone_bd_ram_n19478, 
        p_wishbone_bd_ram_n19479, p_wishbone_bd_ram_n19480, 
        p_wishbone_bd_ram_n19481, p_wishbone_bd_ram_n19482, 
        p_wishbone_bd_ram_n19483, p_wishbone_bd_ram_n19484, 
        p_wishbone_bd_ram_n19485, p_wishbone_bd_ram_n19486, 
        p_wishbone_bd_ram_n19487, p_wishbone_bd_ram_n19488, 
        p_wishbone_bd_ram_n19489, p_wishbone_bd_ram_n19490, 
        p_wishbone_bd_ram_n19491, p_wishbone_bd_ram_n19492, 
        p_wishbone_bd_ram_n19493, p_wishbone_bd_ram_n19494, 
        p_wishbone_bd_ram_n19495, p_wishbone_bd_ram_n19496, 
        p_wishbone_bd_ram_n19497, p_wishbone_bd_ram_n19498, 
        p_wishbone_bd_ram_n19499, p_wishbone_bd_ram_n19500, 
        p_wishbone_bd_ram_n19501, p_wishbone_bd_ram_n19502, 
        p_wishbone_bd_ram_n19503, p_wishbone_bd_ram_n19504, 
        p_wishbone_bd_ram_n19505, p_wishbone_bd_ram_n19506, 
        p_wishbone_bd_ram_n19507, p_wishbone_bd_ram_n19508, 
        p_wishbone_bd_ram_n19509, p_wishbone_bd_ram_n19510, 
        p_wishbone_bd_ram_n19511, p_wishbone_bd_ram_n19512, 
        p_wishbone_bd_ram_n19513, p_wishbone_bd_ram_n19514, 
        p_wishbone_bd_ram_n19515, p_wishbone_bd_ram_n19516, 
        p_wishbone_bd_ram_n19517, p_wishbone_bd_ram_n19518, 
        p_wishbone_bd_ram_n19519, p_wishbone_bd_ram_n19520, 
        p_wishbone_bd_ram_n19521, p_wishbone_bd_ram_n19522, 
        p_wishbone_bd_ram_n19523, p_wishbone_bd_ram_n19524, 
        p_wishbone_bd_ram_n19525, p_wishbone_bd_ram_n19526, 
        p_wishbone_bd_ram_n19527, p_wishbone_bd_ram_n19528, 
        p_wishbone_bd_ram_n19529, p_wishbone_bd_ram_n19530, 
        p_wishbone_bd_ram_n19531, p_wishbone_bd_ram_n19532, 
        p_wishbone_bd_ram_n19533, p_wishbone_bd_ram_n19534, 
        p_wishbone_bd_ram_n19535, p_wishbone_bd_ram_n19536, 
        p_wishbone_bd_ram_n19537, p_wishbone_bd_ram_n19538, 
        p_wishbone_bd_ram_n19539, p_wishbone_bd_ram_n19540, 
        p_wishbone_bd_ram_n19541, p_wishbone_bd_ram_n19542, 
        p_wishbone_bd_ram_n19543, p_wishbone_bd_ram_n19544, 
        p_wishbone_bd_ram_n19545, p_wishbone_bd_ram_n19546, 
        p_wishbone_bd_ram_n19547, p_wishbone_bd_ram_n19548, 
        p_wishbone_bd_ram_n19549, p_wishbone_bd_ram_n19550, 
        p_wishbone_bd_ram_n19551, p_wishbone_bd_ram_n19552, 
        p_wishbone_bd_ram_n19553, p_wishbone_bd_ram_n19554, 
        p_wishbone_bd_ram_n19555, p_wishbone_bd_ram_n19556, 
        p_wishbone_bd_ram_n19557, p_wishbone_bd_ram_n19558, 
        p_wishbone_bd_ram_n19559, p_wishbone_bd_ram_n19560, 
        p_wishbone_bd_ram_n19561, p_wishbone_bd_ram_n19562, 
        p_wishbone_bd_ram_n19563, p_wishbone_bd_ram_n19564, 
        p_wishbone_bd_ram_n19565, p_wishbone_bd_ram_n19566, 
        p_wishbone_bd_ram_n19567, p_wishbone_bd_ram_n19568, 
        p_wishbone_bd_ram_n19569, p_wishbone_bd_ram_n19570, 
        p_wishbone_bd_ram_n19571, p_wishbone_bd_ram_n19572, 
        p_wishbone_bd_ram_n19573, p_wishbone_bd_ram_n19574, 
        p_wishbone_bd_ram_n19575, p_wishbone_bd_ram_n19576, 
        p_wishbone_bd_ram_n19577, p_wishbone_bd_ram_n19578, 
        p_wishbone_bd_ram_n19579, p_wishbone_bd_ram_n19580, 
        p_wishbone_bd_ram_n19581, p_wishbone_bd_ram_n19582, 
        p_wishbone_bd_ram_n19583, p_wishbone_bd_ram_n19584, 
        p_wishbone_bd_ram_n19585, p_wishbone_bd_ram_n19586, 
        p_wishbone_bd_ram_n19587, p_wishbone_bd_ram_n19588, 
        p_wishbone_bd_ram_n19589, p_wishbone_bd_ram_n19590, 
        p_wishbone_bd_ram_n19591, p_wishbone_bd_ram_n19592, 
        p_wishbone_bd_ram_n19593, p_wishbone_bd_ram_n19594, 
        p_wishbone_bd_ram_n19595, p_wishbone_bd_ram_n19596, 
        p_wishbone_bd_ram_n19597, p_wishbone_bd_ram_n19598, 
        p_wishbone_bd_ram_n19599, p_wishbone_bd_ram_n19600, 
        p_wishbone_bd_ram_n19601, p_wishbone_bd_ram_n19602, 
        p_wishbone_bd_ram_n19603, p_wishbone_bd_ram_n19604, 
        p_wishbone_bd_ram_n19605, p_wishbone_bd_ram_n19606, 
        p_wishbone_bd_ram_n19607, p_wishbone_bd_ram_n19608, 
        p_wishbone_bd_ram_n19609, p_wishbone_bd_ram_n19610, 
        p_wishbone_bd_ram_n19611, p_wishbone_bd_ram_n19612, 
        p_wishbone_bd_ram_n19613, p_wishbone_bd_ram_n19614, 
        p_wishbone_bd_ram_n19615, p_wishbone_bd_ram_n19616, 
        p_wishbone_bd_ram_n19617, p_wishbone_bd_ram_n19618, 
        p_wishbone_bd_ram_n19619, p_wishbone_bd_ram_n19620, 
        p_wishbone_bd_ram_n19621, p_wishbone_bd_ram_n19622, 
        p_wishbone_bd_ram_n19623, p_wishbone_bd_ram_n19624, 
        p_wishbone_bd_ram_n19625, p_wishbone_bd_ram_n19626, 
        p_wishbone_bd_ram_n19627, p_wishbone_bd_ram_n19628, 
        p_wishbone_bd_ram_n19629, p_wishbone_bd_ram_n19630, 
        p_wishbone_bd_ram_n19631, p_wishbone_bd_ram_n19632, 
        p_wishbone_bd_ram_n19633, p_wishbone_bd_ram_n19634, 
        p_wishbone_bd_ram_n19635, p_wishbone_bd_ram_n19636, 
        p_wishbone_bd_ram_n19637, p_wishbone_bd_ram_n19638, 
        p_wishbone_bd_ram_n19639, p_wishbone_bd_ram_n19640, 
        p_wishbone_bd_ram_n19641, p_wishbone_bd_ram_n19642, 
        p_wishbone_bd_ram_n19643, p_wishbone_bd_ram_n19644, 
        p_wishbone_bd_ram_n19645, p_wishbone_bd_ram_n19646, 
        p_wishbone_bd_ram_n19647, p_wishbone_bd_ram_n19648, 
        p_wishbone_bd_ram_n19649, p_wishbone_bd_ram_n19650, 
        p_wishbone_bd_ram_n19651, p_wishbone_bd_ram_n19652, 
        p_wishbone_bd_ram_n19653, p_wishbone_bd_ram_n19654, 
        p_wishbone_bd_ram_n19655, p_wishbone_bd_ram_n19656, 
        p_wishbone_bd_ram_n19657, p_wishbone_bd_ram_n19658, 
        p_wishbone_bd_ram_n19659, p_wishbone_bd_ram_n19660, 
        p_wishbone_bd_ram_n19661, p_wishbone_bd_ram_n19662, 
        p_wishbone_bd_ram_n19663, p_wishbone_bd_ram_n19664, 
        p_wishbone_bd_ram_n19665, p_wishbone_bd_ram_n19666, 
        p_wishbone_bd_ram_n19667, p_wishbone_bd_ram_n19668, 
        p_wishbone_bd_ram_n19669, p_wishbone_bd_ram_n19670, 
        p_wishbone_bd_ram_n19671, p_wishbone_bd_ram_n19672, 
        p_wishbone_bd_ram_n19673, p_wishbone_bd_ram_n19674, 
        p_wishbone_bd_ram_n19675, p_wishbone_bd_ram_n19676, 
        p_wishbone_bd_ram_n19677, p_wishbone_bd_ram_n19678, 
        p_wishbone_bd_ram_n19679, p_wishbone_bd_ram_n19680, 
        p_wishbone_bd_ram_n19681, p_wishbone_bd_ram_n19682, 
        p_wishbone_bd_ram_n19683, p_wishbone_bd_ram_n19684, 
        p_wishbone_bd_ram_n19685, p_wishbone_bd_ram_n19686, 
        p_wishbone_bd_ram_n19687, p_wishbone_bd_ram_n19688, 
        p_wishbone_bd_ram_n19689, p_wishbone_bd_ram_n19690, 
        p_wishbone_bd_ram_n19691, p_wishbone_bd_ram_n19692, 
        p_wishbone_bd_ram_n19693, p_wishbone_bd_ram_n19694, 
        p_wishbone_bd_ram_n19695, p_wishbone_bd_ram_n19696, 
        p_wishbone_bd_ram_n19697, p_wishbone_bd_ram_n19698, 
        p_wishbone_bd_ram_n19699, p_wishbone_bd_ram_n19700, 
        p_wishbone_bd_ram_n19701, p_wishbone_bd_ram_n19702, 
        p_wishbone_bd_ram_n19703, p_wishbone_bd_ram_n19704, 
        p_wishbone_bd_ram_n19705, p_wishbone_bd_ram_n19706, 
        p_wishbone_bd_ram_n19707, p_wishbone_bd_ram_n19708, 
        p_wishbone_bd_ram_n19709, p_wishbone_bd_ram_n19710, 
        p_wishbone_bd_ram_n19711, p_wishbone_bd_ram_n19712, 
        p_wishbone_bd_ram_n19713, p_wishbone_bd_ram_n19714, 
        p_wishbone_bd_ram_n19715, p_wishbone_bd_ram_n19716, 
        p_wishbone_bd_ram_n19717, p_wishbone_bd_ram_n19718, 
        p_wishbone_bd_ram_n19719, p_wishbone_bd_ram_n19720, 
        p_wishbone_bd_ram_n19721, p_wishbone_bd_ram_n19722, 
        p_wishbone_bd_ram_n19723, p_wishbone_bd_ram_n19724, 
        p_wishbone_bd_ram_n19725, p_wishbone_bd_ram_n19726, 
        p_wishbone_bd_ram_n19727, p_wishbone_bd_ram_n19728, 
        p_wishbone_bd_ram_n19729, p_wishbone_bd_ram_n19730, 
        p_wishbone_bd_ram_n19731, p_wishbone_bd_ram_n19732, 
        p_wishbone_bd_ram_n19733, p_wishbone_bd_ram_n19734, 
        p_wishbone_bd_ram_n19735, p_wishbone_bd_ram_n19736, 
        p_wishbone_bd_ram_n19737, p_wishbone_bd_ram_n19738, 
        p_wishbone_bd_ram_n19739, p_wishbone_bd_ram_n19740, 
        p_wishbone_bd_ram_n19741, p_wishbone_bd_ram_n19742, 
        p_wishbone_bd_ram_n19743, p_wishbone_bd_ram_n19744, 
        p_wishbone_bd_ram_n19745, p_wishbone_bd_ram_n19746, 
        p_wishbone_bd_ram_n19747, p_wishbone_bd_ram_n19748, 
        p_wishbone_bd_ram_n19749, p_wishbone_bd_ram_n19750, 
        p_wishbone_bd_ram_n19751, p_wishbone_bd_ram_n19752, 
        p_wishbone_bd_ram_n19753, p_wishbone_bd_ram_n19754, 
        p_wishbone_bd_ram_n19755, p_wishbone_bd_ram_n19756, 
        p_wishbone_bd_ram_n19757, p_wishbone_bd_ram_n19758, 
        p_wishbone_bd_ram_n19759, p_wishbone_bd_ram_n19760, 
        p_wishbone_bd_ram_n19761, p_wishbone_bd_ram_n19762, 
        p_wishbone_bd_ram_n19763, p_wishbone_bd_ram_n19764, 
        p_wishbone_bd_ram_n19765, p_wishbone_bd_ram_n19766, 
        p_wishbone_bd_ram_n19767, p_wishbone_bd_ram_n19768, 
        p_wishbone_bd_ram_n19769, p_wishbone_bd_ram_n19770, 
        p_wishbone_bd_ram_n19771, p_wishbone_bd_ram_n19772, 
        p_wishbone_bd_ram_n19773, p_wishbone_bd_ram_n19774, 
        p_wishbone_bd_ram_n19775, p_wishbone_bd_ram_n19776, 
        p_wishbone_bd_ram_n19777, p_wishbone_bd_ram_n19778, 
        p_wishbone_bd_ram_n19779, p_wishbone_bd_ram_n19780, 
        p_wishbone_bd_ram_n19781, p_wishbone_bd_ram_n19782, 
        p_wishbone_bd_ram_n19783, p_wishbone_bd_ram_n19784, 
        p_wishbone_bd_ram_n19785, p_wishbone_bd_ram_n19786, 
        p_wishbone_bd_ram_n19787, p_wishbone_bd_ram_n19788, 
        p_wishbone_bd_ram_n19789, p_wishbone_bd_ram_n19790, 
        p_wishbone_bd_ram_n19791, p_wishbone_bd_ram_n19792, 
        p_wishbone_bd_ram_n19793, p_wishbone_bd_ram_n19794, 
        p_wishbone_bd_ram_n19795, p_wishbone_bd_ram_n19796, 
        p_wishbone_bd_ram_n19797, p_wishbone_bd_ram_n19798, 
        p_wishbone_bd_ram_n19799, p_wishbone_bd_ram_n19800, 
        p_wishbone_bd_ram_n19801, p_wishbone_bd_ram_n19802, 
        p_wishbone_bd_ram_n19803, p_wishbone_bd_ram_n19804, 
        p_wishbone_bd_ram_n19805, p_wishbone_bd_ram_n19806, 
        p_wishbone_bd_ram_n19807, p_wishbone_bd_ram_n19808, 
        p_wishbone_bd_ram_n19809, p_wishbone_bd_ram_n19810, 
        p_wishbone_bd_ram_n19811, p_wishbone_bd_ram_n19812, 
        p_wishbone_bd_ram_n19813, p_wishbone_bd_ram_n19814, 
        p_wishbone_bd_ram_n19815, p_wishbone_bd_ram_n19816, 
        p_wishbone_bd_ram_n19817, p_wishbone_bd_ram_n19818, 
        p_wishbone_bd_ram_n19819, p_wishbone_bd_ram_n19820, 
        p_wishbone_bd_ram_n19821, p_wishbone_bd_ram_n19822, 
        p_wishbone_bd_ram_n19823, p_wishbone_bd_ram_n19824, 
        p_wishbone_bd_ram_n19825, p_wishbone_bd_ram_n19826, 
        p_wishbone_bd_ram_n19827, p_wishbone_bd_ram_n19828, 
        p_wishbone_bd_ram_n19829, p_wishbone_bd_ram_n19830, 
        p_wishbone_bd_ram_n19831, p_wishbone_bd_ram_n19832, 
        p_wishbone_bd_ram_n19833, p_wishbone_bd_ram_n19834, 
        p_wishbone_bd_ram_n19835, p_wishbone_bd_ram_n19836, 
        p_wishbone_bd_ram_n19837, p_wishbone_bd_ram_n19838, 
        p_wishbone_bd_ram_n19839, p_wishbone_bd_ram_n19840, 
        p_wishbone_bd_ram_n19841, p_wishbone_bd_ram_n19842, 
        p_wishbone_bd_ram_n19843, p_wishbone_bd_ram_n19844, 
        p_wishbone_bd_ram_n19845, p_wishbone_bd_ram_n19846, 
        p_wishbone_bd_ram_n19847, p_wishbone_bd_ram_n19848, 
        p_wishbone_bd_ram_n19849, p_wishbone_bd_ram_n19850, 
        p_wishbone_bd_ram_n19851, p_wishbone_bd_ram_n19852, 
        p_wishbone_bd_ram_n19853, p_wishbone_bd_ram_n19854, 
        p_wishbone_bd_ram_n19855, p_wishbone_bd_ram_n19856, 
        p_wishbone_bd_ram_n19857, p_wishbone_bd_ram_n19858, 
        p_wishbone_bd_ram_n19859, p_wishbone_bd_ram_n19860, 
        p_wishbone_bd_ram_n19861, p_wishbone_bd_ram_n19862, 
        p_wishbone_bd_ram_n19863, p_wishbone_bd_ram_n19864, 
        p_wishbone_bd_ram_n19865, p_wishbone_bd_ram_n19866, 
        p_wishbone_bd_ram_n19867, p_wishbone_bd_ram_n19868, 
        p_wishbone_bd_ram_n19869, p_wishbone_bd_ram_n19870, 
        p_wishbone_bd_ram_n19871, p_wishbone_bd_ram_n19872, 
        p_wishbone_bd_ram_n19873, p_wishbone_bd_ram_n19874, 
        p_wishbone_bd_ram_n19875, p_wishbone_bd_ram_n19876, 
        p_wishbone_bd_ram_n19877, p_wishbone_bd_ram_n19878, 
        p_wishbone_bd_ram_n19879, p_wishbone_bd_ram_n19880, 
        p_wishbone_bd_ram_n19881, p_wishbone_bd_ram_n19882, 
        p_wishbone_bd_ram_n19883, p_wishbone_bd_ram_n19884, 
        p_wishbone_bd_ram_n19885, p_wishbone_bd_ram_n19886, 
        p_wishbone_bd_ram_n19887, p_wishbone_bd_ram_n19888, 
        p_wishbone_bd_ram_n19889, p_wishbone_bd_ram_n19890, 
        p_wishbone_bd_ram_n19891, p_wishbone_bd_ram_n19892, 
        p_wishbone_bd_ram_n19893, p_wishbone_bd_ram_n19894, 
        p_wishbone_bd_ram_n19895, p_wishbone_bd_ram_n19896, 
        p_wishbone_bd_ram_n19897, p_wishbone_bd_ram_n19898, 
        p_wishbone_bd_ram_n19899, p_wishbone_bd_ram_n19900, 
        p_wishbone_bd_ram_n19901, p_wishbone_bd_ram_n19902, 
        p_wishbone_bd_ram_n19903, p_wishbone_bd_ram_n19904, 
        p_wishbone_bd_ram_n19905, p_wishbone_bd_ram_n19906, 
        p_wishbone_bd_ram_n19907, p_wishbone_bd_ram_n19908, 
        p_wishbone_bd_ram_n19909, p_wishbone_bd_ram_n19910, 
        p_wishbone_bd_ram_n19911, p_wishbone_bd_ram_n19912, 
        p_wishbone_bd_ram_n19913, p_wishbone_bd_ram_n19914, 
        p_wishbone_bd_ram_n19915, p_wishbone_bd_ram_n19916, 
        p_wishbone_bd_ram_n19917, p_wishbone_bd_ram_n19918, 
        p_wishbone_bd_ram_n19919, p_wishbone_bd_ram_n19920, 
        p_wishbone_bd_ram_n19921, p_wishbone_bd_ram_n19922, 
        p_wishbone_bd_ram_n19923, p_wishbone_bd_ram_n19924, 
        p_wishbone_bd_ram_n19925, p_wishbone_bd_ram_n19926, 
        p_wishbone_bd_ram_n19927, p_wishbone_bd_ram_n19928, 
        p_wishbone_bd_ram_n19929, p_wishbone_bd_ram_n19930, 
        p_wishbone_bd_ram_n19931, p_wishbone_bd_ram_n19932, 
        p_wishbone_bd_ram_n19933, p_wishbone_bd_ram_n19934, 
        p_wishbone_bd_ram_n19935, p_wishbone_bd_ram_n19936, 
        p_wishbone_bd_ram_n19937, p_wishbone_bd_ram_n19938, 
        p_wishbone_bd_ram_n19939, p_wishbone_bd_ram_n19940, 
        p_wishbone_bd_ram_n19941, p_wishbone_bd_ram_n19942, 
        p_wishbone_bd_ram_n19943, p_wishbone_bd_ram_n19944, 
        p_wishbone_bd_ram_n19945, p_wishbone_bd_ram_n19946, 
        p_wishbone_bd_ram_n19947, p_wishbone_bd_ram_n19948, 
        p_wishbone_bd_ram_n19949, p_wishbone_bd_ram_n19950, 
        p_wishbone_bd_ram_n19951, p_wishbone_bd_ram_n19952, 
        p_wishbone_bd_ram_n19953, p_wishbone_bd_ram_n19954, 
        p_wishbone_bd_ram_n19955, p_wishbone_bd_ram_n19956, 
        p_wishbone_bd_ram_n19957, p_wishbone_bd_ram_n19958, 
        p_wishbone_bd_ram_n19959, p_wishbone_bd_ram_n19960, 
        p_wishbone_bd_ram_n19961, p_wishbone_bd_ram_n19962, 
        p_wishbone_bd_ram_n19963, p_wishbone_bd_ram_n19964, 
        p_wishbone_bd_ram_n19965, p_wishbone_bd_ram_n19966, 
        p_wishbone_bd_ram_n19967, p_wishbone_bd_ram_n19968, 
        p_wishbone_bd_ram_n19969, p_wishbone_bd_ram_n19970, 
        p_wishbone_bd_ram_n19971, p_wishbone_bd_ram_n19972, 
        p_wishbone_bd_ram_n19973, p_wishbone_bd_ram_n19974, 
        p_wishbone_bd_ram_n19975, p_wishbone_bd_ram_n19976, 
        p_wishbone_bd_ram_n19977, p_wishbone_bd_ram_n19978, 
        p_wishbone_bd_ram_n19979, p_wishbone_bd_ram_n19980, 
        p_wishbone_bd_ram_n19981, p_wishbone_bd_ram_n19982, 
        p_wishbone_bd_ram_n19983, p_wishbone_bd_ram_n19984, 
        p_wishbone_bd_ram_n19985, p_wishbone_bd_ram_n19986, 
        p_wishbone_bd_ram_n19987, p_wishbone_bd_ram_n19988, 
        p_wishbone_bd_ram_n19989, p_wishbone_bd_ram_n19990, 
        p_wishbone_bd_ram_n19991, p_wishbone_bd_ram_n19992, 
        p_wishbone_bd_ram_n19993, p_wishbone_bd_ram_n19994, 
        p_wishbone_bd_ram_n19995, p_wishbone_bd_ram_n19996, 
        p_wishbone_bd_ram_n19997, p_wishbone_bd_ram_n19998, 
        p_wishbone_bd_ram_n19999, p_wishbone_bd_ram_n20000, 
        p_wishbone_bd_ram_n20001, p_wishbone_bd_ram_n20002, 
        p_wishbone_bd_ram_n20003, p_wishbone_bd_ram_n20004, 
        p_wishbone_bd_ram_n20005, p_wishbone_bd_ram_n20006, 
        p_wishbone_bd_ram_n20007, p_wishbone_bd_ram_n20008, 
        p_wishbone_bd_ram_n20009, p_wishbone_bd_ram_n20010, 
        p_wishbone_bd_ram_n20011, p_wishbone_bd_ram_n20012, 
        p_wishbone_bd_ram_n20013, p_wishbone_bd_ram_n20014, 
        p_wishbone_bd_ram_n20015, p_wishbone_bd_ram_n20016, 
        p_wishbone_bd_ram_n20017, p_wishbone_bd_ram_n20018, 
        p_wishbone_bd_ram_n20019, p_wishbone_bd_ram_n20020, 
        p_wishbone_bd_ram_n20021, p_wishbone_bd_ram_n20022, 
        p_wishbone_bd_ram_n20023, p_wishbone_bd_ram_n20024, 
        p_wishbone_bd_ram_n20025, p_wishbone_bd_ram_n20026, 
        p_wishbone_bd_ram_n20027, p_wishbone_bd_ram_n20028, 
        p_wishbone_bd_ram_n20029, p_wishbone_bd_ram_n20030, 
        p_wishbone_bd_ram_n20031, p_wishbone_bd_ram_n20032, 
        p_wishbone_bd_ram_n20033, p_wishbone_bd_ram_n20034, 
        p_wishbone_bd_ram_n20035, p_wishbone_bd_ram_n20036, 
        p_wishbone_bd_ram_n20037, p_wishbone_bd_ram_n20038, 
        p_wishbone_bd_ram_n20039, p_wishbone_bd_ram_n20040, 
        p_wishbone_bd_ram_n20041, p_wishbone_bd_ram_n20042, 
        p_wishbone_bd_ram_n20043, p_wishbone_bd_ram_n20044, 
        p_wishbone_bd_ram_n20045, p_wishbone_bd_ram_n20046, 
        p_wishbone_bd_ram_n20047, p_wishbone_bd_ram_n20048, 
        p_wishbone_bd_ram_n20049, p_wishbone_bd_ram_n20050, 
        p_wishbone_bd_ram_n20051, p_wishbone_bd_ram_n20052, 
        p_wishbone_bd_ram_n20053, p_wishbone_bd_ram_n20054, 
        p_wishbone_bd_ram_n20055, p_wishbone_bd_ram_n20056, 
        p_wishbone_bd_ram_n20057, p_wishbone_bd_ram_n20058, 
        p_wishbone_bd_ram_n20059, p_wishbone_bd_ram_n20060, 
        p_wishbone_bd_ram_n20061, p_wishbone_bd_ram_n20062, 
        p_wishbone_bd_ram_n20063, p_wishbone_bd_ram_n20064, 
        p_wishbone_bd_ram_n20065, p_wishbone_bd_ram_n20066, 
        p_wishbone_bd_ram_n20067, p_wishbone_bd_ram_n20068, 
        p_wishbone_bd_ram_n20069, p_wishbone_bd_ram_n20070, 
        p_wishbone_bd_ram_n20071, p_wishbone_bd_ram_n20072, 
        p_wishbone_bd_ram_n20073, p_wishbone_bd_ram_n20074, 
        p_wishbone_bd_ram_n20075, p_wishbone_bd_ram_n20076, 
        p_wishbone_bd_ram_n20077, p_wishbone_bd_ram_n20078, 
        p_wishbone_bd_ram_n20079, p_wishbone_bd_ram_n20080, 
        p_wishbone_bd_ram_n20081, p_wishbone_bd_ram_n20082, 
        p_wishbone_bd_ram_n20083, p_wishbone_bd_ram_n20084, 
        p_wishbone_bd_ram_n20085, p_wishbone_bd_ram_n20086, 
        p_wishbone_bd_ram_n20087, p_wishbone_bd_ram_n20088, 
        p_wishbone_bd_ram_n20089, p_wishbone_bd_ram_n20090, 
        p_wishbone_bd_ram_n20091, p_wishbone_bd_ram_n20092, 
        p_wishbone_bd_ram_n20093, p_wishbone_bd_ram_n20094, 
        p_wishbone_bd_ram_n20095, p_wishbone_bd_ram_n20096, 
        p_wishbone_bd_ram_n20097, p_wishbone_bd_ram_n20098, 
        p_wishbone_bd_ram_n20099, p_wishbone_bd_ram_n20100, 
        p_wishbone_bd_ram_n20101, p_wishbone_bd_ram_n20102, 
        p_wishbone_bd_ram_n20103, p_wishbone_bd_ram_n20104, 
        p_wishbone_bd_ram_n20105, p_wishbone_bd_ram_n20106, 
        p_wishbone_bd_ram_n20107, p_wishbone_bd_ram_n20108, 
        p_wishbone_bd_ram_n20109, p_wishbone_bd_ram_n20110, 
        p_wishbone_bd_ram_n20111, p_wishbone_bd_ram_n20112, 
        p_wishbone_bd_ram_n20113, p_wishbone_bd_ram_n20114, 
        p_wishbone_bd_ram_n20115, p_wishbone_bd_ram_n20116, 
        p_wishbone_bd_ram_n20117, p_wishbone_bd_ram_n20118, 
        p_wishbone_bd_ram_n20119, p_wishbone_bd_ram_n20120, 
        p_wishbone_bd_ram_n20121, p_wishbone_bd_ram_n20122, 
        p_wishbone_bd_ram_n20123, p_wishbone_bd_ram_n20124, 
        p_wishbone_bd_ram_n20125, p_wishbone_bd_ram_n20126, 
        p_wishbone_bd_ram_n20127, p_wishbone_bd_ram_n20128, 
        p_wishbone_bd_ram_n20129, p_wishbone_bd_ram_n20130, 
        p_wishbone_bd_ram_n20131, p_wishbone_bd_ram_n20132, 
        p_wishbone_bd_ram_n20133, p_wishbone_bd_ram_n20134, 
        p_wishbone_bd_ram_n20135, p_wishbone_bd_ram_n20136, 
        p_wishbone_bd_ram_n20137, p_wishbone_bd_ram_n20138, 
        p_wishbone_bd_ram_n20139, p_wishbone_bd_ram_n20140, 
        p_wishbone_bd_ram_n20141, p_wishbone_bd_ram_n20142, 
        p_wishbone_bd_ram_n20143, p_wishbone_bd_ram_n20144, 
        p_wishbone_bd_ram_n20145, p_wishbone_bd_ram_n20146, 
        p_wishbone_bd_ram_n20147, p_wishbone_bd_ram_n20148, 
        p_wishbone_bd_ram_n20149, p_wishbone_bd_ram_n20150, 
        p_wishbone_bd_ram_n20151, p_wishbone_bd_ram_n20152, 
        p_wishbone_bd_ram_n20153, p_wishbone_bd_ram_n20154, 
        p_wishbone_bd_ram_n20155, p_wishbone_bd_ram_n20156, 
        p_wishbone_bd_ram_n20157, p_wishbone_bd_ram_n20158, 
        p_wishbone_bd_ram_n20159, p_wishbone_bd_ram_n20160, 
        p_wishbone_bd_ram_n20161, p_wishbone_bd_ram_n20162, 
        p_wishbone_bd_ram_n20163, p_wishbone_bd_ram_n20164, 
        p_wishbone_bd_ram_n20165, p_wishbone_bd_ram_n20166, 
        p_wishbone_bd_ram_n20167, p_wishbone_bd_ram_n20168, 
        p_wishbone_bd_ram_n20169, p_wishbone_bd_ram_n20170, 
        p_wishbone_bd_ram_n20171, p_wishbone_bd_ram_n20172, 
        p_wishbone_bd_ram_n20173, p_wishbone_bd_ram_n20174, 
        p_wishbone_bd_ram_n20175, p_wishbone_bd_ram_n20176, 
        p_wishbone_bd_ram_n20177, p_wishbone_bd_ram_n20178, 
        p_wishbone_bd_ram_n20179, p_wishbone_bd_ram_n20180, 
        p_wishbone_bd_ram_n20181, p_wishbone_bd_ram_n20182, 
        p_wishbone_bd_ram_n20183, p_wishbone_bd_ram_n20184, 
        p_wishbone_bd_ram_n20185, p_wishbone_bd_ram_n20186, 
        p_wishbone_bd_ram_n20187, p_wishbone_bd_ram_n20188, 
        p_wishbone_bd_ram_n20189, p_wishbone_bd_ram_n20190, 
        p_wishbone_bd_ram_n20191, p_wishbone_bd_ram_n20192, 
        p_wishbone_bd_ram_n20193, p_wishbone_bd_ram_n20194, 
        p_wishbone_bd_ram_n20195, p_wishbone_bd_ram_n20196, 
        p_wishbone_bd_ram_n20197, p_wishbone_bd_ram_n20198, 
        p_wishbone_bd_ram_n20199, p_wishbone_bd_ram_n20200, 
        p_wishbone_bd_ram_n20201, p_wishbone_bd_ram_n20202, 
        p_wishbone_bd_ram_n20203, p_wishbone_bd_ram_n20204, 
        p_wishbone_bd_ram_n20205, p_wishbone_bd_ram_n20206, 
        p_wishbone_bd_ram_n20207, p_wishbone_bd_ram_n20208, 
        p_wishbone_bd_ram_n20209, p_wishbone_bd_ram_n20210, 
        p_wishbone_bd_ram_n20211, p_wishbone_bd_ram_n20212, 
        p_wishbone_bd_ram_n20213, p_wishbone_bd_ram_n20214, 
        p_wishbone_bd_ram_n20215, p_wishbone_bd_ram_n20216, 
        p_wishbone_bd_ram_n20217, p_wishbone_bd_ram_n20218, 
        p_wishbone_bd_ram_n20219, p_wishbone_bd_ram_n20220, 
        p_wishbone_bd_ram_n20221, p_wishbone_bd_ram_n20222, 
        p_wishbone_bd_ram_n20223, p_wishbone_bd_ram_n20224, 
        p_wishbone_bd_ram_n20225, p_wishbone_bd_ram_n20226, 
        p_wishbone_bd_ram_n20227, p_wishbone_bd_ram_n20228, 
        p_wishbone_bd_ram_n20229, p_wishbone_bd_ram_n20230, 
        p_wishbone_bd_ram_n20231, p_wishbone_bd_ram_n20232, 
        p_wishbone_bd_ram_n20233, p_wishbone_bd_ram_n20234, 
        p_wishbone_bd_ram_n20235, p_wishbone_bd_ram_n20236, 
        p_wishbone_bd_ram_n20237, p_wishbone_bd_ram_n20238, 
        p_wishbone_bd_ram_n20239, p_wishbone_bd_ram_n20240, 
        p_wishbone_bd_ram_n20241, p_wishbone_bd_ram_n20242, 
        p_wishbone_bd_ram_n20243, p_wishbone_bd_ram_n20244, 
        p_wishbone_bd_ram_n20245, p_wishbone_bd_ram_n20246, 
        p_wishbone_bd_ram_n20247, p_wishbone_bd_ram_n20248, 
        p_wishbone_bd_ram_n20249, p_wishbone_bd_ram_n20250, 
        p_wishbone_bd_ram_n20251, p_wishbone_bd_ram_n20252, 
        p_wishbone_bd_ram_n20253, p_wishbone_bd_ram_n20254, 
        p_wishbone_bd_ram_n20255, p_wishbone_bd_ram_n20256, 
        p_wishbone_bd_ram_n20257, p_wishbone_bd_ram_n20258, 
        p_wishbone_bd_ram_n20259, p_wishbone_bd_ram_n20260, 
        p_wishbone_bd_ram_n20261, p_wishbone_bd_ram_n20262, 
        p_wishbone_bd_ram_n20263, p_wishbone_bd_ram_n20264, 
        p_wishbone_bd_ram_n20265, p_wishbone_bd_ram_n20266, 
        p_wishbone_bd_ram_n20267, p_wishbone_bd_ram_n20268, 
        p_wishbone_bd_ram_n20269, p_wishbone_bd_ram_n20270, 
        p_wishbone_bd_ram_n20271, p_wishbone_bd_ram_n20272, 
        p_wishbone_bd_ram_n20273, p_wishbone_bd_ram_n20274, 
        p_wishbone_bd_ram_n20275, p_wishbone_bd_ram_n20276, 
        p_wishbone_bd_ram_n20277, p_wishbone_bd_ram_n20278, 
        p_wishbone_bd_ram_n20279, p_wishbone_bd_ram_n20280, 
        p_wishbone_bd_ram_n20281, p_wishbone_bd_ram_n20282, 
        p_wishbone_bd_ram_n20283, p_wishbone_bd_ram_n20284, 
        p_wishbone_bd_ram_n20285, p_wishbone_bd_ram_n20286, 
        p_wishbone_bd_ram_n20287, p_wishbone_bd_ram_n20288, 
        p_wishbone_bd_ram_n20289, p_wishbone_bd_ram_n20290, 
        p_wishbone_bd_ram_n20291, p_wishbone_bd_ram_n20292, 
        p_wishbone_bd_ram_n20293, p_wishbone_bd_ram_n20294, 
        p_wishbone_bd_ram_n20295, p_wishbone_bd_ram_n20296, 
        p_wishbone_bd_ram_n20297, p_wishbone_bd_ram_n20298, 
        p_wishbone_bd_ram_n20299, p_wishbone_bd_ram_n20300, 
        p_wishbone_bd_ram_n20301, p_wishbone_bd_ram_n20302, 
        p_wishbone_bd_ram_n20303, p_wishbone_bd_ram_n20304, 
        p_wishbone_bd_ram_n20305, p_wishbone_bd_ram_n20306, 
        p_wishbone_bd_ram_n20307, p_wishbone_bd_ram_n20308, 
        p_wishbone_bd_ram_n20309, p_wishbone_bd_ram_n20310, 
        p_wishbone_bd_ram_n20311, p_wishbone_bd_ram_n20312, 
        p_wishbone_bd_ram_n20313, p_wishbone_bd_ram_n20314, 
        p_wishbone_bd_ram_n20315, p_wishbone_bd_ram_n20316, 
        p_wishbone_bd_ram_n20317, p_wishbone_bd_ram_n20318, 
        p_wishbone_bd_ram_n20319, p_wishbone_bd_ram_n20320, 
        p_wishbone_bd_ram_n20321, p_wishbone_bd_ram_n20322, 
        p_wishbone_bd_ram_n20323, p_wishbone_bd_ram_n20324, 
        p_wishbone_bd_ram_n20325, p_wishbone_bd_ram_n20326, 
        p_wishbone_bd_ram_n20327, p_wishbone_bd_ram_n20328, 
        p_wishbone_bd_ram_n20329, p_wishbone_bd_ram_n20330, 
        p_wishbone_bd_ram_n20331, p_wishbone_bd_ram_n20332, 
        p_wishbone_bd_ram_n20333, p_wishbone_bd_ram_n20334, 
        p_wishbone_bd_ram_n20335, p_wishbone_bd_ram_n20336, 
        p_wishbone_bd_ram_n20337, p_wishbone_bd_ram_n20338, 
        p_wishbone_bd_ram_n20339, p_wishbone_bd_ram_n20340, 
        p_wishbone_bd_ram_n20341, p_wishbone_bd_ram_n20342, 
        p_wishbone_bd_ram_n20343, p_wishbone_bd_ram_n20344, 
        p_wishbone_bd_ram_n20345, p_wishbone_bd_ram_n20346, 
        p_wishbone_bd_ram_n20347, p_wishbone_bd_ram_n20348, 
        p_wishbone_bd_ram_n20349, p_wishbone_bd_ram_n20350, 
        p_wishbone_bd_ram_n20351, p_wishbone_bd_ram_n20352, 
        p_wishbone_bd_ram_n20353, p_wishbone_bd_ram_n20354, 
        p_wishbone_bd_ram_n20355, p_wishbone_bd_ram_n20356, 
        p_wishbone_bd_ram_n20357, p_wishbone_bd_ram_n20358, 
        p_wishbone_bd_ram_n20359, p_wishbone_bd_ram_n20360, 
        p_wishbone_bd_ram_n20361, p_wishbone_bd_ram_n20362, 
        p_wishbone_bd_ram_n20363, p_wishbone_bd_ram_n20364, 
        p_wishbone_bd_ram_n20365, p_wishbone_bd_ram_n20366, 
        p_wishbone_bd_ram_n20367, p_wishbone_bd_ram_n20368, 
        p_wishbone_bd_ram_n20369, p_wishbone_bd_ram_n20370, 
        p_wishbone_bd_ram_n20371, p_wishbone_bd_ram_n20372, 
        p_wishbone_bd_ram_n20373, p_wishbone_bd_ram_n20374, 
        p_wishbone_bd_ram_n20375, p_wishbone_bd_ram_n20376, 
        p_wishbone_bd_ram_n20377, p_wishbone_bd_ram_n20378, 
        p_wishbone_bd_ram_n20379, p_wishbone_bd_ram_n20380, 
        p_wishbone_bd_ram_n20381, p_wishbone_bd_ram_n20382, 
        p_wishbone_bd_ram_n20383, p_wishbone_bd_ram_n20384, 
        p_wishbone_bd_ram_n20385, p_wishbone_bd_ram_n20386, 
        p_wishbone_bd_ram_n20387, p_wishbone_bd_ram_n20388, 
        p_wishbone_bd_ram_n20389, p_wishbone_bd_ram_n20390, 
        p_wishbone_bd_ram_n20391, p_wishbone_bd_ram_n20392, 
        p_wishbone_bd_ram_n20393, p_wishbone_bd_ram_n20394, 
        p_wishbone_bd_ram_n20395, p_wishbone_bd_ram_n20396, 
        p_wishbone_bd_ram_n20397, p_wishbone_bd_ram_n20398, 
        p_wishbone_bd_ram_n20399, p_wishbone_bd_ram_n20400, 
        p_wishbone_bd_ram_n20401, p_wishbone_bd_ram_n20402, 
        p_wishbone_bd_ram_n20403, p_wishbone_bd_ram_n20404, 
        p_wishbone_bd_ram_n20405, p_wishbone_bd_ram_n20406, 
        p_wishbone_bd_ram_n20407, p_wishbone_bd_ram_n20408, 
        p_wishbone_bd_ram_n20409, p_wishbone_bd_ram_n20410, 
        p_wishbone_bd_ram_n20411, p_wishbone_bd_ram_n20412, 
        p_wishbone_bd_ram_n20413, p_wishbone_bd_ram_n20414, 
        p_wishbone_bd_ram_n20415, p_wishbone_bd_ram_n20416, 
        p_wishbone_bd_ram_n20417, p_wishbone_bd_ram_n20418, 
        p_wishbone_bd_ram_n20419, p_wishbone_bd_ram_n20420, 
        p_wishbone_bd_ram_n20421, p_wishbone_bd_ram_n20422, 
        p_wishbone_bd_ram_n20423, p_wishbone_bd_ram_n20424, 
        p_wishbone_bd_ram_n20425, p_wishbone_bd_ram_n20426, 
        p_wishbone_bd_ram_n20427, p_wishbone_bd_ram_n20428, 
        p_wishbone_bd_ram_n20429, p_wishbone_bd_ram_n20430, 
        p_wishbone_bd_ram_n20431, p_wishbone_bd_ram_n20432, 
        p_wishbone_bd_ram_n20433, p_wishbone_bd_ram_n20434, 
        p_wishbone_bd_ram_n20435, p_wishbone_bd_ram_n20436, 
        p_wishbone_bd_ram_n20437, p_wishbone_bd_ram_n20438, 
        p_wishbone_bd_ram_n20439, p_wishbone_bd_ram_n20440, 
        p_wishbone_bd_ram_n20441, p_wishbone_bd_ram_n20442, 
        p_wishbone_bd_ram_n20443, p_wishbone_bd_ram_n20444, 
        p_wishbone_bd_ram_n20445, p_wishbone_bd_ram_n20446, 
        p_wishbone_bd_ram_n20447, p_wishbone_bd_ram_n20448, 
        p_wishbone_bd_ram_n20449, p_wishbone_bd_ram_n20450, 
        p_wishbone_bd_ram_n20451, p_wishbone_bd_ram_n20452, 
        p_wishbone_bd_ram_n20453, p_wishbone_bd_ram_n20454, 
        p_wishbone_bd_ram_n20455, p_wishbone_bd_ram_n20456, 
        p_wishbone_bd_ram_n20457, p_wishbone_bd_ram_n20458, 
        p_wishbone_bd_ram_n20459, p_wishbone_bd_ram_n20460, 
        p_wishbone_bd_ram_n20461, p_wishbone_bd_ram_n20462, 
        p_wishbone_bd_ram_n20463, p_wishbone_bd_ram_n20464, 
        p_wishbone_bd_ram_n20465, p_wishbone_bd_ram_n20466, 
        p_wishbone_bd_ram_n20467, p_wishbone_bd_ram_n20468, 
        p_wishbone_bd_ram_n20469, p_wishbone_bd_ram_n20470, 
        p_wishbone_bd_ram_n20471, p_wishbone_bd_ram_n20472, 
        p_wishbone_bd_ram_n20473, p_wishbone_bd_ram_n20474, 
        p_wishbone_bd_ram_n20475, p_wishbone_bd_ram_n20476, 
        p_wishbone_bd_ram_n20477, p_wishbone_bd_ram_n20478, 
        p_wishbone_bd_ram_n20479, p_wishbone_bd_ram_n20480, 
        p_wishbone_bd_ram_n20481, p_wishbone_bd_ram_n20482, 
        p_wishbone_bd_ram_n20483, p_wishbone_bd_ram_n20484, 
        p_wishbone_bd_ram_n20485, p_wishbone_bd_ram_n20486, 
        p_wishbone_bd_ram_n20487, p_wishbone_bd_ram_n20488, 
        p_wishbone_bd_ram_n20489, p_wishbone_bd_ram_n20490, 
        p_wishbone_bd_ram_n20491, p_wishbone_bd_ram_n20492, 
        p_wishbone_bd_ram_n20493, p_wishbone_bd_ram_n20494, 
        p_wishbone_bd_ram_n20495, p_wishbone_bd_ram_n20496, 
        p_wishbone_bd_ram_n20497, p_wishbone_bd_ram_n20498, 
        p_wishbone_bd_ram_n20499, p_wishbone_bd_ram_n20500, 
        p_wishbone_bd_ram_n20501, p_wishbone_bd_ram_n20502, 
        p_wishbone_bd_ram_n20503, p_wishbone_bd_ram_n20504, 
        p_wishbone_bd_ram_n20505, p_wishbone_bd_ram_n20506, 
        p_wishbone_bd_ram_n20507, p_wishbone_bd_ram_n20508, 
        p_wishbone_bd_ram_n20509, p_wishbone_bd_ram_n20510, 
        p_wishbone_bd_ram_n20511, p_wishbone_bd_ram_n20512, 
        p_wishbone_bd_ram_n20513, p_wishbone_bd_ram_n20514, 
        p_wishbone_bd_ram_n20515, p_wishbone_bd_ram_n20516, 
        p_wishbone_bd_ram_n20517, p_wishbone_bd_ram_n20518, 
        p_wishbone_bd_ram_n20519, p_wishbone_bd_ram_n20520, 
        p_wishbone_bd_ram_n20521, p_wishbone_bd_ram_n20522, 
        p_wishbone_bd_ram_n20523, p_wishbone_bd_ram_n20524, 
        p_wishbone_bd_ram_n20525, p_wishbone_bd_ram_n20526, 
        p_wishbone_bd_ram_n20527, p_wishbone_bd_ram_n20528, 
        p_wishbone_bd_ram_n20529, p_wishbone_bd_ram_n20530, 
        p_wishbone_bd_ram_n20531, p_wishbone_bd_ram_n20532, 
        p_wishbone_bd_ram_n20533, p_wishbone_bd_ram_n20534, 
        p_wishbone_bd_ram_n20535, p_wishbone_bd_ram_n20536, 
        p_wishbone_bd_ram_n20537, p_wishbone_bd_ram_n20538, 
        p_wishbone_bd_ram_n20539, p_wishbone_bd_ram_n20540, 
        p_wishbone_bd_ram_n20541, p_wishbone_bd_ram_n20542, 
        p_wishbone_bd_ram_n20543, p_wishbone_bd_ram_n20544, 
        p_wishbone_bd_ram_n20545, p_wishbone_bd_ram_n20546, 
        p_wishbone_bd_ram_n20547, p_wishbone_bd_ram_n20548, 
        p_wishbone_bd_ram_n20549, p_wishbone_bd_ram_n20550, 
        p_wishbone_bd_ram_n20551, p_wishbone_bd_ram_n20552, 
        p_wishbone_bd_ram_n20553, p_wishbone_bd_ram_n20554, 
        p_wishbone_bd_ram_n20555, p_wishbone_bd_ram_n20556, 
        p_wishbone_bd_ram_n20557, p_wishbone_bd_ram_n20558, 
        p_wishbone_bd_ram_n20559, p_wishbone_bd_ram_n20560, 
        p_wishbone_bd_ram_n20561, p_wishbone_bd_ram_n20562, 
        p_wishbone_bd_ram_n20563, p_wishbone_bd_ram_n20564, 
        p_wishbone_bd_ram_n20565, p_wishbone_bd_ram_n20566, 
        p_wishbone_bd_ram_n20567, p_wishbone_bd_ram_n20568, 
        p_wishbone_bd_ram_n20569, p_wishbone_bd_ram_n20570, 
        p_wishbone_bd_ram_n20571, p_wishbone_bd_ram_n20572, 
        p_wishbone_bd_ram_n20573, p_wishbone_bd_ram_n20574, 
        p_wishbone_bd_ram_n20575, p_wishbone_bd_ram_n20576, 
        p_wishbone_bd_ram_n20577, p_wishbone_bd_ram_n20578, 
        p_wishbone_bd_ram_n20579, p_wishbone_bd_ram_n20580, 
        p_wishbone_bd_ram_n20581, p_wishbone_bd_ram_n20582, 
        p_wishbone_bd_ram_n20583, p_wishbone_bd_ram_n20584, 
        p_wishbone_bd_ram_n20585, p_wishbone_bd_ram_n20586, 
        p_wishbone_bd_ram_n20587, p_wishbone_bd_ram_n20588, 
        p_wishbone_bd_ram_n20589, p_wishbone_bd_ram_n20590, 
        p_wishbone_bd_ram_n20591, p_wishbone_bd_ram_n20592, 
        p_wishbone_bd_ram_n20593, p_wishbone_bd_ram_n20594, 
        p_wishbone_bd_ram_n20595, p_wishbone_bd_ram_n20596, 
        p_wishbone_bd_ram_n20597, p_wishbone_bd_ram_n20598, 
        p_wishbone_bd_ram_n20599, p_wishbone_bd_ram_n20600, 
        p_wishbone_bd_ram_n20601, p_wishbone_bd_ram_n20602, 
        p_wishbone_bd_ram_n20603, p_wishbone_bd_ram_n20604, 
        p_wishbone_bd_ram_n20605, p_wishbone_bd_ram_n20606, 
        p_wishbone_bd_ram_n20607, p_wishbone_bd_ram_n20608, 
        p_wishbone_bd_ram_n20609, p_wishbone_bd_ram_n20610, 
        p_wishbone_bd_ram_n20611, p_wishbone_bd_ram_n20612, 
        p_wishbone_bd_ram_n20613, p_wishbone_bd_ram_n20614, 
        p_wishbone_bd_ram_n20615, p_wishbone_bd_ram_n20616, 
        p_wishbone_bd_ram_n20617, p_wishbone_bd_ram_n20618, 
        p_wishbone_bd_ram_n20619, p_wishbone_bd_ram_n20620, 
        p_wishbone_bd_ram_n20621, p_wishbone_bd_ram_n20622, 
        p_wishbone_bd_ram_n20623, p_wishbone_bd_ram_n20624, 
        p_wishbone_bd_ram_n20625, p_wishbone_bd_ram_n20626, 
        p_wishbone_bd_ram_n20627, p_wishbone_bd_ram_n20628, 
        p_wishbone_bd_ram_n20629, p_wishbone_bd_ram_n20630, 
        p_wishbone_bd_ram_n20631, p_wishbone_bd_ram_n20632, 
        p_wishbone_bd_ram_n20633, p_wishbone_bd_ram_n20634, 
        p_wishbone_bd_ram_n20635, p_wishbone_bd_ram_n20636, 
        p_wishbone_bd_ram_n20637, p_wishbone_bd_ram_n20638, 
        p_wishbone_bd_ram_n20639, p_wishbone_bd_ram_n20640, 
        p_wishbone_bd_ram_n20641, p_wishbone_bd_ram_n20642, 
        p_wishbone_bd_ram_n20643, p_wishbone_bd_ram_n20644, 
        p_wishbone_bd_ram_n20645, p_wishbone_bd_ram_n20646, 
        p_wishbone_bd_ram_n20647, p_wishbone_bd_ram_n20648, 
        p_wishbone_bd_ram_n20649, p_wishbone_bd_ram_n20650, 
        p_wishbone_bd_ram_n20651, p_wishbone_bd_ram_n20652, 
        p_wishbone_bd_ram_n20653, p_wishbone_bd_ram_n20654, 
        p_wishbone_bd_ram_n20655, p_wishbone_bd_ram_n20656, 
        p_wishbone_bd_ram_n20657, p_wishbone_bd_ram_n20658, 
        p_wishbone_bd_ram_n20659, p_wishbone_bd_ram_n20660, 
        p_wishbone_bd_ram_n20661, p_wishbone_bd_ram_n20662, 
        p_wishbone_bd_ram_n20663, p_wishbone_bd_ram_n20664, 
        p_wishbone_bd_ram_n20665, p_wishbone_bd_ram_n20666, 
        p_wishbone_bd_ram_n20667, p_wishbone_bd_ram_n20668, 
        p_wishbone_bd_ram_n20669, p_wishbone_bd_ram_n20670, 
        p_wishbone_bd_ram_n20671, p_wishbone_bd_ram_n20672, 
        p_wishbone_bd_ram_n20673, p_wishbone_bd_ram_n20674, 
        p_wishbone_bd_ram_n20675, p_wishbone_bd_ram_n20676, 
        p_wishbone_bd_ram_n20677, p_wishbone_bd_ram_n20678, 
        p_wishbone_bd_ram_n20679, p_wishbone_bd_ram_n20680, 
        p_wishbone_bd_ram_n20681, p_wishbone_bd_ram_n20682, 
        p_wishbone_bd_ram_n20683, p_wishbone_bd_ram_n20684, 
        p_wishbone_bd_ram_n20685, p_wishbone_bd_ram_n20686, 
        p_wishbone_bd_ram_n20687, p_wishbone_bd_ram_n20688, 
        p_wishbone_bd_ram_n20689, p_wishbone_bd_ram_n20690, 
        p_wishbone_bd_ram_n20691, p_wishbone_bd_ram_n20692, 
        p_wishbone_bd_ram_n20693, p_wishbone_bd_ram_n20694, 
        p_wishbone_bd_ram_n20695, p_wishbone_bd_ram_n20696, 
        p_wishbone_bd_ram_n20697, p_wishbone_bd_ram_n20698, 
        p_wishbone_bd_ram_n20699, p_wishbone_bd_ram_n20700, 
        p_wishbone_bd_ram_n20701, p_wishbone_bd_ram_n20702, 
        p_wishbone_bd_ram_n20703, p_wishbone_bd_ram_n20704, 
        p_wishbone_bd_ram_n20705, p_wishbone_bd_ram_n20706, 
        p_wishbone_bd_ram_n20707, p_wishbone_bd_ram_n20708, 
        p_wishbone_bd_ram_n20709, p_wishbone_bd_ram_n20710, 
        p_wishbone_bd_ram_n20711, p_wishbone_bd_ram_n20712, 
        p_wishbone_bd_ram_n20713, p_wishbone_bd_ram_n20714, 
        p_wishbone_bd_ram_n20715, p_wishbone_bd_ram_n20716, 
        p_wishbone_bd_ram_n20717, p_wishbone_bd_ram_n20718, 
        p_wishbone_bd_ram_n20719, p_wishbone_bd_ram_n20720, 
        p_wishbone_bd_ram_n20721, p_wishbone_bd_ram_n20722, 
        p_wishbone_bd_ram_n20723, p_wishbone_bd_ram_n20724, 
        p_wishbone_bd_ram_n20725, p_wishbone_bd_ram_n20726, 
        p_wishbone_bd_ram_n20727, p_wishbone_bd_ram_n20728, 
        p_wishbone_bd_ram_n20729, p_wishbone_bd_ram_n20730, 
        p_wishbone_bd_ram_n20731, p_wishbone_bd_ram_n20732, 
        p_wishbone_bd_ram_n20733, p_wishbone_bd_ram_n20734, 
        p_wishbone_bd_ram_n20735, p_wishbone_bd_ram_n20736, 
        p_wishbone_bd_ram_n20737, p_wishbone_bd_ram_n20738, 
        p_wishbone_bd_ram_n20739, p_wishbone_bd_ram_n20740, 
        p_wishbone_bd_ram_n20741, p_wishbone_bd_ram_n20742, 
        p_wishbone_bd_ram_n20743, p_wishbone_bd_ram_n20744, 
        p_wishbone_bd_ram_n20745, p_wishbone_bd_ram_n20746, 
        p_wishbone_bd_ram_n20747, p_wishbone_bd_ram_n20748, 
        p_wishbone_bd_ram_n20749, p_wishbone_bd_ram_n20750, 
        p_wishbone_bd_ram_n20751, p_wishbone_bd_ram_n20752, 
        p_wishbone_bd_ram_n20753, p_wishbone_bd_ram_n20754, 
        p_wishbone_bd_ram_n20755, p_wishbone_bd_ram_n20756, 
        p_wishbone_bd_ram_n20757, p_wishbone_bd_ram_n20758, 
        p_wishbone_bd_ram_n20759, p_wishbone_bd_ram_n20760, 
        p_wishbone_bd_ram_n20761, p_wishbone_bd_ram_n20762, 
        p_wishbone_bd_ram_n20763, p_wishbone_bd_ram_n20764, 
        p_wishbone_bd_ram_n20765, p_wishbone_bd_ram_n20766, 
        p_wishbone_bd_ram_n20767, p_wishbone_bd_ram_n20768, 
        p_wishbone_bd_ram_n20769, p_wishbone_bd_ram_n20770, 
        p_wishbone_bd_ram_n20771, p_wishbone_bd_ram_n20772, 
        p_wishbone_bd_ram_n20773, p_wishbone_bd_ram_n20774, 
        p_wishbone_bd_ram_n20775, p_wishbone_bd_ram_n20776, 
        p_wishbone_bd_ram_n20777, p_wishbone_bd_ram_n20778, 
        p_wishbone_bd_ram_n20779, p_wishbone_bd_ram_n20780, 
        p_wishbone_bd_ram_n20781, p_wishbone_bd_ram_n20782, 
        p_wishbone_bd_ram_n20783, p_wishbone_bd_ram_n20784, 
        p_wishbone_bd_ram_n20785, p_wishbone_bd_ram_n20786, 
        p_wishbone_bd_ram_n20787, p_wishbone_bd_ram_n20788, 
        p_wishbone_bd_ram_n20789, p_wishbone_bd_ram_n20790, 
        p_wishbone_bd_ram_n20791, p_wishbone_bd_ram_n20792, 
        p_wishbone_bd_ram_n20793, p_wishbone_bd_ram_n20794, 
        p_wishbone_bd_ram_n20795, p_wishbone_bd_ram_n20796, 
        p_wishbone_bd_ram_n20797, p_wishbone_bd_ram_n20798, 
        p_wishbone_bd_ram_n20799, p_wishbone_bd_ram_n20800, 
        p_wishbone_bd_ram_n20801, p_wishbone_bd_ram_n20802, 
        p_wishbone_bd_ram_n20803, p_wishbone_bd_ram_n20804, 
        p_wishbone_bd_ram_n20805, p_wishbone_bd_ram_n20806, 
        p_wishbone_bd_ram_n20807, p_wishbone_bd_ram_n20808, 
        p_wishbone_bd_ram_n20809, p_wishbone_bd_ram_n20810, 
        p_wishbone_bd_ram_n20811, p_wishbone_bd_ram_n20812, 
        p_wishbone_bd_ram_n20813, p_wishbone_bd_ram_n20814, 
        p_wishbone_bd_ram_n20815, p_wishbone_bd_ram_n20816, 
        p_wishbone_bd_ram_n20817, p_wishbone_bd_ram_n20818, 
        p_wishbone_bd_ram_n20819, p_wishbone_bd_ram_n20820, 
        p_wishbone_bd_ram_n20821, p_wishbone_bd_ram_n20822, 
        p_wishbone_bd_ram_n20823, p_wishbone_bd_ram_n20824, 
        p_wishbone_bd_ram_n20825, p_wishbone_bd_ram_n20826, 
        p_wishbone_bd_ram_n20827, p_wishbone_bd_ram_n20828, 
        p_wishbone_bd_ram_n20829, p_wishbone_bd_ram_n20830, 
        p_wishbone_bd_ram_n20831, p_wishbone_bd_ram_n20832, 
        p_wishbone_bd_ram_n20833, p_wishbone_bd_ram_n20834, 
        p_wishbone_bd_ram_n20835, p_wishbone_bd_ram_n20836, 
        p_wishbone_bd_ram_n20837, p_wishbone_bd_ram_n20838, 
        p_wishbone_bd_ram_n20839, p_wishbone_bd_ram_n20840, 
        p_wishbone_bd_ram_n20841, p_wishbone_bd_ram_n20842, 
        p_wishbone_bd_ram_n20843, p_wishbone_bd_ram_n20844, 
        p_wishbone_bd_ram_n20845, p_wishbone_bd_ram_n20846, 
        p_wishbone_bd_ram_n20847, p_wishbone_bd_ram_n20848, 
        p_wishbone_bd_ram_n20849, p_wishbone_bd_ram_n20850, 
        p_wishbone_bd_ram_n20851, p_wishbone_bd_ram_n20852, 
        p_wishbone_bd_ram_n20853, p_wishbone_bd_ram_n20854, 
        p_wishbone_bd_ram_n20855, p_wishbone_bd_ram_n20856, 
        p_wishbone_bd_ram_n20857, p_wishbone_bd_ram_n20858, 
        p_wishbone_bd_ram_n20859, p_wishbone_bd_ram_n20860, 
        p_wishbone_bd_ram_n20861, p_wishbone_bd_ram_n20862, 
        p_wishbone_bd_ram_n20863, p_wishbone_bd_ram_n20864, 
        p_wishbone_bd_ram_n20865, p_wishbone_bd_ram_n20866, 
        p_wishbone_bd_ram_n20867, p_wishbone_bd_ram_n20868, 
        p_wishbone_bd_ram_n20869, p_wishbone_bd_ram_n20870, 
        p_wishbone_bd_ram_n20871, p_wishbone_bd_ram_n20872, 
        p_wishbone_bd_ram_n20873, p_wishbone_bd_ram_n20874, 
        p_wishbone_bd_ram_n20875, p_wishbone_bd_ram_n20876, 
        p_wishbone_bd_ram_n20877, p_wishbone_bd_ram_n20878, 
        p_wishbone_bd_ram_n20879, p_wishbone_bd_ram_n20880, 
        p_wishbone_bd_ram_n20881, p_wishbone_bd_ram_n20882, 
        p_wishbone_bd_ram_n20883, p_wishbone_bd_ram_n20884, 
        p_wishbone_bd_ram_n20885, p_wishbone_bd_ram_n20886, 
        p_wishbone_bd_ram_n20887, p_wishbone_bd_ram_n20888, 
        p_wishbone_bd_ram_n20889, p_wishbone_bd_ram_n20890, 
        p_wishbone_bd_ram_n20891, p_wishbone_bd_ram_n20892, 
        p_wishbone_bd_ram_n20893, p_wishbone_bd_ram_n20894, 
        p_wishbone_bd_ram_n20895, p_wishbone_bd_ram_n20896, 
        p_wishbone_bd_ram_n20897, p_wishbone_bd_ram_n20898, 
        p_wishbone_bd_ram_n20899, p_wishbone_bd_ram_n20900, 
        p_wishbone_bd_ram_n20901, p_wishbone_bd_ram_n20902, 
        p_wishbone_bd_ram_n20903, p_wishbone_bd_ram_n20904, 
        p_wishbone_bd_ram_n20905, p_wishbone_bd_ram_n20906, 
        p_wishbone_bd_ram_n20907, p_wishbone_bd_ram_n20908, 
        p_wishbone_bd_ram_n20909, p_wishbone_bd_ram_n20910, 
        p_wishbone_bd_ram_n20911, p_wishbone_bd_ram_n20912, 
        p_wishbone_bd_ram_n20913, p_wishbone_bd_ram_n20914, 
        p_wishbone_bd_ram_n20915, p_wishbone_bd_ram_n20916, 
        p_wishbone_bd_ram_n20917, p_wishbone_bd_ram_n20918, 
        p_wishbone_bd_ram_n20919, p_wishbone_bd_ram_n20920, 
        p_wishbone_bd_ram_n20921, p_wishbone_bd_ram_n20922, 
        p_wishbone_bd_ram_n20923, p_wishbone_bd_ram_n20924, 
        p_wishbone_bd_ram_n20925, p_wishbone_bd_ram_n20926, 
        p_wishbone_bd_ram_n20927, p_wishbone_bd_ram_n20928, 
        p_wishbone_bd_ram_n20929, p_wishbone_bd_ram_n20930, 
        p_wishbone_bd_ram_n20931, p_wishbone_bd_ram_n20932, 
        p_wishbone_bd_ram_n20933, p_wishbone_bd_ram_n20934, 
        p_wishbone_bd_ram_n20935, p_wishbone_bd_ram_n20936, 
        p_wishbone_bd_ram_n20937, p_wishbone_bd_ram_n20938, 
        p_wishbone_bd_ram_n20939, p_wishbone_bd_ram_n20940, 
        p_wishbone_bd_ram_n20941, p_wishbone_bd_ram_n20942, 
        p_wishbone_bd_ram_n20943, p_wishbone_bd_ram_n20944, 
        p_wishbone_bd_ram_n20945, p_wishbone_bd_ram_n20946, 
        p_wishbone_bd_ram_n20947, p_wishbone_bd_ram_n20948, 
        p_wishbone_bd_ram_n20949, p_wishbone_bd_ram_n20950, 
        p_wishbone_bd_ram_n20951, p_wishbone_bd_ram_n20952, 
        p_wishbone_bd_ram_n20953, p_wishbone_bd_ram_n20954, 
        p_wishbone_bd_ram_n20955, p_wishbone_bd_ram_n20956, 
        p_wishbone_bd_ram_n20957, p_wishbone_bd_ram_n20958, 
        p_wishbone_bd_ram_n20959, p_wishbone_bd_ram_n20960, 
        p_wishbone_bd_ram_n20961, p_wishbone_bd_ram_n20962, 
        p_wishbone_bd_ram_n20963, p_wishbone_bd_ram_n20964, 
        p_wishbone_bd_ram_n20965, p_wishbone_bd_ram_n20966, 
        p_wishbone_bd_ram_n20967, p_wishbone_bd_ram_n20968, 
        p_wishbone_bd_ram_n20969, p_wishbone_bd_ram_n20970, 
        p_wishbone_bd_ram_n20971, p_wishbone_bd_ram_n20972, 
        p_wishbone_bd_ram_n20973, p_wishbone_bd_ram_n20974, 
        p_wishbone_bd_ram_n20975, p_wishbone_bd_ram_n20976, 
        p_wishbone_bd_ram_n20977, p_wishbone_bd_ram_n20978, 
        p_wishbone_bd_ram_n20979, p_wishbone_bd_ram_n20980, 
        p_wishbone_bd_ram_n20981, p_wishbone_bd_ram_n20982, 
        p_wishbone_bd_ram_n20983, p_wishbone_bd_ram_n20984, 
        p_wishbone_bd_ram_n20985, p_wishbone_bd_ram_n20986, 
        p_wishbone_bd_ram_n20987, p_wishbone_bd_ram_n20988, 
        p_wishbone_bd_ram_n20989, p_wishbone_bd_ram_n20990, 
        p_wishbone_bd_ram_n20991, p_wishbone_bd_ram_n20992, 
        p_wishbone_bd_ram_n20993, p_wishbone_bd_ram_n20994, 
        p_wishbone_bd_ram_n20995, p_wishbone_bd_ram_n20996, 
        p_wishbone_bd_ram_n20997, p_wishbone_bd_ram_n20998, 
        p_wishbone_bd_ram_n20999, p_wishbone_bd_ram_n21000, 
        p_wishbone_bd_ram_n21001, p_wishbone_bd_ram_n21002, 
        p_wishbone_bd_ram_n21003, p_wishbone_bd_ram_n21004, 
        p_wishbone_bd_ram_n21005, p_wishbone_bd_ram_n21006, 
        p_wishbone_bd_ram_n21007, p_wishbone_bd_ram_n21008, 
        p_wishbone_bd_ram_n21009, p_wishbone_bd_ram_n21010, 
        p_wishbone_bd_ram_n21011, p_wishbone_bd_ram_n21012, 
        p_wishbone_bd_ram_n21013, p_wishbone_bd_ram_n21014, 
        p_wishbone_bd_ram_n21015, p_wishbone_bd_ram_n21016, 
        p_wishbone_bd_ram_n21017, p_wishbone_bd_ram_n21018, 
        p_wishbone_bd_ram_n21019, p_wishbone_bd_ram_n21020, 
        p_wishbone_bd_ram_n21021, p_wishbone_bd_ram_n21022, 
        p_wishbone_bd_ram_n21023, p_wishbone_bd_ram_n21024, 
        p_wishbone_bd_ram_n21025, p_wishbone_bd_ram_n21026, 
        p_wishbone_bd_ram_n21027, p_wishbone_bd_ram_n21028, 
        p_wishbone_bd_ram_n21029, p_wishbone_bd_ram_n21030, 
        p_wishbone_bd_ram_n21031, p_wishbone_bd_ram_n21032, 
        p_wishbone_bd_ram_n21033, p_wishbone_bd_ram_n21034, 
        p_wishbone_bd_ram_n21035, p_wishbone_bd_ram_n21036, 
        p_wishbone_bd_ram_n21037, p_wishbone_bd_ram_n21038, 
        p_wishbone_bd_ram_n21039, p_wishbone_bd_ram_n21040, 
        p_wishbone_bd_ram_n21041, p_wishbone_bd_ram_n21042, 
        p_wishbone_bd_ram_n21043, p_wishbone_bd_ram_n21044, 
        p_wishbone_bd_ram_n21045, p_wishbone_bd_ram_n21046, 
        p_wishbone_bd_ram_n21047, p_wishbone_bd_ram_n21048, 
        p_wishbone_bd_ram_n21049, p_wishbone_bd_ram_n21050, 
        p_wishbone_bd_ram_n21051, p_wishbone_bd_ram_n21052, 
        p_wishbone_bd_ram_n21053, p_wishbone_bd_ram_n21054, 
        p_wishbone_bd_ram_n21055, p_wishbone_bd_ram_n21056, 
        p_wishbone_bd_ram_n21057, p_wishbone_bd_ram_n21058, 
        p_wishbone_bd_ram_n21059, p_wishbone_bd_ram_n21060, 
        p_wishbone_bd_ram_n21061, p_wishbone_bd_ram_n21062, 
        p_wishbone_bd_ram_n21063, p_wishbone_bd_ram_n21064, 
        p_wishbone_bd_ram_n21065, p_wishbone_bd_ram_n21066, 
        p_wishbone_bd_ram_n21067, p_wishbone_bd_ram_n21068, 
        p_wishbone_bd_ram_n21069, p_wishbone_bd_ram_n21070, 
        p_wishbone_bd_ram_n21071, p_wishbone_bd_ram_n21072, 
        p_wishbone_bd_ram_n21073, p_wishbone_bd_ram_n21074, 
        p_wishbone_bd_ram_n21075, p_wishbone_bd_ram_n21076, 
        p_wishbone_bd_ram_n21077, p_wishbone_bd_ram_n21078, 
        p_wishbone_bd_ram_n21079, p_wishbone_bd_ram_n21080, 
        p_wishbone_bd_ram_n21081, p_wishbone_bd_ram_n21082, 
        p_wishbone_bd_ram_n21083, p_wishbone_bd_ram_n21084, 
        p_wishbone_bd_ram_n21085, p_wishbone_bd_ram_n21086, 
        p_wishbone_bd_ram_n21087, p_wishbone_bd_ram_n21088, 
        p_wishbone_bd_ram_n21089, p_wishbone_bd_ram_n21090, 
        p_wishbone_bd_ram_n21091, p_wishbone_bd_ram_n21092, 
        p_wishbone_bd_ram_n21093, p_wishbone_bd_ram_n21094, 
        p_wishbone_bd_ram_n21095, p_wishbone_bd_ram_n21096, 
        p_wishbone_bd_ram_n21097, p_wishbone_bd_ram_n21098, 
        p_wishbone_bd_ram_n21099, p_wishbone_bd_ram_n21100, 
        p_wishbone_bd_ram_n21101, p_wishbone_bd_ram_n21102, 
        p_wishbone_bd_ram_n21103, p_wishbone_bd_ram_n21104, 
        p_wishbone_bd_ram_n21105, p_wishbone_bd_ram_n21106, 
        p_wishbone_bd_ram_n21107, p_wishbone_bd_ram_n21108, 
        p_wishbone_bd_ram_n21109, p_wishbone_bd_ram_n21110, 
        p_wishbone_bd_ram_n21111, p_wishbone_bd_ram_n21112, 
        p_wishbone_bd_ram_n21113, p_wishbone_bd_ram_n21114, 
        p_wishbone_bd_ram_n21115, p_wishbone_bd_ram_n21116, 
        p_wishbone_bd_ram_n21117, p_wishbone_bd_ram_n21118, 
        p_wishbone_bd_ram_n21119, p_wishbone_bd_ram_n21120, 
        p_wishbone_bd_ram_n21121, p_wishbone_bd_ram_n21122, 
        p_wishbone_bd_ram_n21123, p_wishbone_bd_ram_n21124, 
        p_wishbone_bd_ram_n21125, p_wishbone_bd_ram_n21126, 
        p_wishbone_bd_ram_n21127, p_wishbone_bd_ram_n21128, 
        p_wishbone_bd_ram_n21129, p_wishbone_bd_ram_n21130, 
        p_wishbone_bd_ram_n21131, p_wishbone_bd_ram_n21132, 
        p_wishbone_bd_ram_n21133, p_wishbone_bd_ram_n21134, 
        p_wishbone_bd_ram_n21135, p_wishbone_bd_ram_n21136, 
        p_wishbone_bd_ram_n21137, p_wishbone_bd_ram_n21138, 
        p_wishbone_bd_ram_n21139, p_wishbone_bd_ram_n21140, 
        p_wishbone_bd_ram_n21141, p_wishbone_bd_ram_n21142, 
        p_wishbone_bd_ram_n21143, p_wishbone_bd_ram_n21144, 
        p_wishbone_bd_ram_n21145, p_wishbone_bd_ram_n21146, 
        p_wishbone_bd_ram_n21147, p_wishbone_bd_ram_n21148, 
        p_wishbone_bd_ram_n21149, p_wishbone_bd_ram_n21150, 
        p_wishbone_bd_ram_n21151, p_wishbone_bd_ram_n21152, 
        p_wishbone_bd_ram_n21153, p_wishbone_bd_ram_n21154, 
        p_wishbone_bd_ram_n21155, p_wishbone_bd_ram_n21156, 
        p_wishbone_bd_ram_n21157, p_wishbone_bd_ram_n21158, 
        p_wishbone_bd_ram_n21159, p_wishbone_bd_ram_n21160, 
        p_wishbone_bd_ram_n21161, p_wishbone_bd_ram_n21162, 
        p_wishbone_bd_ram_n21163, p_wishbone_bd_ram_n21164, 
        p_wishbone_bd_ram_n21165, p_wishbone_bd_ram_n21166, 
        p_wishbone_bd_ram_n21167, p_wishbone_bd_ram_n21168, 
        p_wishbone_bd_ram_n21169, p_wishbone_bd_ram_n21170, 
        p_wishbone_bd_ram_n21171, p_wishbone_bd_ram_n21172, 
        p_wishbone_bd_ram_n21173, p_wishbone_bd_ram_n21174, 
        p_wishbone_bd_ram_n21175, p_wishbone_bd_ram_n21176, 
        p_wishbone_bd_ram_n21177, p_wishbone_bd_ram_n21178, 
        p_wishbone_bd_ram_n21179, p_wishbone_bd_ram_n21180, 
        p_wishbone_bd_ram_n21181, p_wishbone_bd_ram_n21182, 
        p_wishbone_bd_ram_n21183, p_wishbone_bd_ram_n21184, 
        p_wishbone_bd_ram_n21185, p_wishbone_bd_ram_n21186, 
        p_wishbone_bd_ram_n21187, p_wishbone_bd_ram_n21188, 
        p_wishbone_bd_ram_n21189, p_wishbone_bd_ram_n21190, 
        p_wishbone_bd_ram_n21191, p_wishbone_bd_ram_n21192, 
        p_wishbone_bd_ram_n21193, p_wishbone_bd_ram_n21194, 
        p_wishbone_bd_ram_n21195, p_wishbone_bd_ram_n21196, 
        p_wishbone_bd_ram_n21197, p_wishbone_bd_ram_n21198, 
        p_wishbone_bd_ram_n21199, p_wishbone_bd_ram_n21200, 
        p_wishbone_bd_ram_n21201, p_wishbone_bd_ram_n21202, 
        p_wishbone_bd_ram_n21203, p_wishbone_bd_ram_n21204, 
        p_wishbone_bd_ram_n21205, p_wishbone_bd_ram_n21206, 
        p_wishbone_bd_ram_n21207, p_wishbone_bd_ram_n21208, 
        p_wishbone_bd_ram_n21209, p_wishbone_bd_ram_n21210, 
        p_wishbone_bd_ram_n21211, p_wishbone_bd_ram_n21212, 
        p_wishbone_bd_ram_n21213, p_wishbone_bd_ram_n21214, 
        p_wishbone_bd_ram_n21215, p_wishbone_bd_ram_n21216, 
        p_wishbone_bd_ram_n21217, p_wishbone_bd_ram_n21218, 
        p_wishbone_bd_ram_n21219, p_wishbone_bd_ram_n21220, 
        p_wishbone_bd_ram_n21221, p_wishbone_bd_ram_n21222, 
        p_wishbone_bd_ram_n21223, p_wishbone_bd_ram_n21224, 
        p_wishbone_bd_ram_n21225, p_wishbone_bd_ram_n21226, 
        p_wishbone_bd_ram_n21227, p_wishbone_bd_ram_n21228, 
        p_wishbone_bd_ram_n21229, p_wishbone_bd_ram_n21230, 
        p_wishbone_bd_ram_n21231, p_wishbone_bd_ram_n21232, 
        p_wishbone_bd_ram_n21233, p_wishbone_bd_ram_n21234, 
        p_wishbone_bd_ram_n21235, p_wishbone_bd_ram_n21236, 
        p_wishbone_bd_ram_n21237, p_wishbone_bd_ram_n21238, 
        p_wishbone_bd_ram_n21239, p_wishbone_bd_ram_n21240, 
        p_wishbone_bd_ram_n21241, p_wishbone_bd_ram_n21242, 
        p_wishbone_bd_ram_n21243, p_wishbone_bd_ram_n21244, 
        p_wishbone_bd_ram_n21245, p_wishbone_bd_ram_n21246, 
        p_wishbone_bd_ram_n21247, p_wishbone_bd_ram_n21248, 
        p_wishbone_bd_ram_n21249, p_wishbone_bd_ram_n21250, 
        p_wishbone_bd_ram_n21251, p_wishbone_bd_ram_n21252, 
        p_wishbone_bd_ram_n21253, p_wishbone_bd_ram_n21254, 
        p_wishbone_bd_ram_n21255, p_wishbone_bd_ram_n21256, 
        p_wishbone_bd_ram_n21257, p_wishbone_bd_ram_n21258, 
        p_wishbone_bd_ram_n21259, p_wishbone_bd_ram_n21260, 
        p_wishbone_bd_ram_n21261, p_wishbone_bd_ram_n21262, 
        p_wishbone_bd_ram_n21263, p_wishbone_bd_ram_n21264, 
        p_wishbone_bd_ram_n21265, p_wishbone_bd_ram_n21266, 
        p_wishbone_bd_ram_n21267, p_wishbone_bd_ram_n21268, 
        p_wishbone_bd_ram_n21269, p_wishbone_bd_ram_n21270, 
        p_wishbone_bd_ram_n21271, p_wishbone_bd_ram_n21272, 
        p_wishbone_bd_ram_n21273, p_wishbone_bd_ram_n21274, 
        p_wishbone_bd_ram_n21275, p_wishbone_bd_ram_n21276, 
        p_wishbone_bd_ram_n21277, p_wishbone_bd_ram_n21278, 
        p_wishbone_bd_ram_n21279, p_wishbone_bd_ram_n21280, 
        p_wishbone_bd_ram_n21281, p_wishbone_bd_ram_n21282, 
        p_wishbone_bd_ram_n21283, p_wishbone_bd_ram_n21284, 
        p_wishbone_bd_ram_n21285, p_wishbone_bd_ram_n21286, 
        p_wishbone_bd_ram_n21287, p_wishbone_bd_ram_n21288, 
        p_wishbone_bd_ram_n21289, p_wishbone_bd_ram_n21290, 
        p_wishbone_bd_ram_n21291, p_wishbone_bd_ram_n21292, 
        p_wishbone_bd_ram_n21293, p_wishbone_bd_ram_n21294, 
        p_wishbone_bd_ram_n21295, p_wishbone_bd_ram_n21296, 
        p_wishbone_bd_ram_n21297, p_wishbone_bd_ram_n21298, 
        p_wishbone_bd_ram_n21299, p_wishbone_bd_ram_n21300, 
        p_wishbone_bd_ram_n21301, p_wishbone_bd_ram_n21302, 
        p_wishbone_bd_ram_n21303, p_wishbone_bd_ram_n21304, 
        p_wishbone_bd_ram_n21305, p_wishbone_bd_ram_n21306, 
        p_wishbone_bd_ram_n21307, p_wishbone_bd_ram_n21308, 
        p_wishbone_bd_ram_n21309, p_wishbone_bd_ram_n21310, 
        p_wishbone_bd_ram_n21311, p_wishbone_bd_ram_n21312, 
        p_wishbone_bd_ram_n21313, p_wishbone_bd_ram_n21314, 
        p_wishbone_bd_ram_n21315, p_wishbone_bd_ram_n21316, 
        p_wishbone_bd_ram_n21317, p_wishbone_bd_ram_n21318, 
        p_wishbone_bd_ram_n21319, p_wishbone_bd_ram_n21320, 
        p_wishbone_bd_ram_n21321, p_wishbone_bd_ram_n21322, 
        p_wishbone_bd_ram_n21323, p_wishbone_bd_ram_n21324, 
        p_wishbone_bd_ram_n21325, p_wishbone_bd_ram_n21326, 
        p_wishbone_bd_ram_n21327, p_wishbone_bd_ram_n21328, 
        p_wishbone_bd_ram_n21329, p_wishbone_bd_ram_n21330, 
        p_wishbone_bd_ram_n21331, p_wishbone_bd_ram_n21332, 
        p_wishbone_bd_ram_n21333, p_wishbone_bd_ram_n21334, 
        p_wishbone_bd_ram_n21335, p_wishbone_bd_ram_n21336, 
        p_wishbone_bd_ram_n21337, p_wishbone_bd_ram_n21338, 
        p_wishbone_bd_ram_n21339, p_wishbone_bd_ram_n21340, 
        p_wishbone_bd_ram_n21341, p_wishbone_bd_ram_n21342, 
        p_wishbone_bd_ram_n21343, p_wishbone_bd_ram_n21344, 
        p_wishbone_bd_ram_n21345, p_wishbone_bd_ram_n21346, 
        p_wishbone_bd_ram_n21347, p_wishbone_bd_ram_n21348, 
        p_wishbone_bd_ram_n21349, p_wishbone_bd_ram_n21350, 
        p_wishbone_bd_ram_n21351, p_wishbone_bd_ram_n21352, 
        p_wishbone_bd_ram_n21353, p_wishbone_bd_ram_n21354, 
        p_wishbone_bd_ram_n21355, p_wishbone_bd_ram_n21356, 
        p_wishbone_bd_ram_n21357, p_wishbone_bd_ram_n21358, 
        p_wishbone_bd_ram_n21359, p_wishbone_bd_ram_n21360, 
        p_wishbone_bd_ram_n21361, p_wishbone_bd_ram_n21362, 
        p_wishbone_bd_ram_n21363, p_wishbone_bd_ram_n21364, 
        p_wishbone_bd_ram_n21365, p_wishbone_bd_ram_n21366, 
        p_wishbone_bd_ram_n21367, p_wishbone_bd_ram_n21368, 
        p_wishbone_bd_ram_n21369, p_wishbone_bd_ram_n21370, 
        p_wishbone_bd_ram_n21371, p_wishbone_bd_ram_n21372, 
        p_wishbone_bd_ram_n21373, p_wishbone_bd_ram_n21374, 
        p_wishbone_bd_ram_n21375, p_wishbone_bd_ram_n21376, 
        p_wishbone_bd_ram_n21377, p_wishbone_bd_ram_n21378, 
        p_wishbone_bd_ram_n21379, p_wishbone_bd_ram_n21380, 
        p_wishbone_bd_ram_n21381, p_wishbone_bd_ram_n21382, 
        p_wishbone_bd_ram_n21383, p_wishbone_bd_ram_n21384, 
        p_wishbone_bd_ram_n21385, p_wishbone_bd_ram_n21386, 
        p_wishbone_bd_ram_n21387, p_wishbone_bd_ram_n21388, 
        p_wishbone_bd_ram_n21389, p_wishbone_bd_ram_n21390, 
        p_wishbone_bd_ram_n21391, p_wishbone_bd_ram_n21392, 
        p_wishbone_bd_ram_n21393, p_wishbone_bd_ram_n21394, 
        p_wishbone_bd_ram_n21395, p_wishbone_bd_ram_n21396, 
        p_wishbone_bd_ram_n21397, p_wishbone_bd_ram_n21398, 
        p_wishbone_bd_ram_n21399, p_wishbone_bd_ram_n21400, 
        p_wishbone_bd_ram_n21401, p_wishbone_bd_ram_n21402, 
        p_wishbone_bd_ram_n21403, p_wishbone_bd_ram_n21404, 
        p_wishbone_bd_ram_n21405, p_wishbone_bd_ram_n21406, 
        p_wishbone_bd_ram_n21407, p_wishbone_bd_ram_n21408, 
        p_wishbone_bd_ram_n21409, p_wishbone_bd_ram_n21410, 
        p_wishbone_bd_ram_n21411, p_wishbone_bd_ram_n21412, 
        p_wishbone_bd_ram_n21413, p_wishbone_bd_ram_n21414, 
        p_wishbone_bd_ram_n21415, p_wishbone_bd_ram_n21416, 
        p_wishbone_bd_ram_n21417, p_wishbone_bd_ram_n21418, 
        p_wishbone_bd_ram_n21419, p_wishbone_bd_ram_n21420, 
        p_wishbone_bd_ram_n21421, p_wishbone_bd_ram_n21422, 
        p_wishbone_bd_ram_n21423, p_wishbone_bd_ram_n21424, 
        p_wishbone_bd_ram_n21425, p_wishbone_bd_ram_n21426, 
        p_wishbone_bd_ram_n21427, p_wishbone_bd_ram_n21428, 
        p_wishbone_bd_ram_n21429, p_wishbone_bd_ram_n21430, 
        p_wishbone_bd_ram_n21431, p_wishbone_bd_ram_n21432, 
        p_wishbone_bd_ram_n21433, p_wishbone_bd_ram_n21434, 
        p_wishbone_bd_ram_n21435, p_wishbone_bd_ram_n21436, 
        p_wishbone_bd_ram_n21437, p_wishbone_bd_ram_n21438, 
        p_wishbone_bd_ram_n21439, p_wishbone_bd_ram_n21440, 
        p_wishbone_bd_ram_n21441, p_wishbone_bd_ram_n21442, 
        p_wishbone_bd_ram_n21443, p_wishbone_bd_ram_n21444, 
        p_wishbone_bd_ram_n21445, p_wishbone_bd_ram_n21446, 
        p_wishbone_bd_ram_n21447, p_wishbone_bd_ram_n21448, 
        p_wishbone_bd_ram_n21449, p_wishbone_bd_ram_n21450, 
        p_wishbone_bd_ram_n21451, p_wishbone_bd_ram_n21452, 
        p_wishbone_bd_ram_n21453, p_wishbone_bd_ram_n21454, 
        p_wishbone_bd_ram_n21455, p_wishbone_bd_ram_n21456, 
        p_wishbone_bd_ram_n21457, p_wishbone_bd_ram_n21458, 
        p_wishbone_bd_ram_n21459, p_wishbone_bd_ram_n21460, 
        p_wishbone_bd_ram_n21461, p_wishbone_bd_ram_n21462, 
        p_wishbone_bd_ram_n21463, p_wishbone_bd_ram_n21464, 
        p_wishbone_bd_ram_n21465, p_wishbone_bd_ram_n21466, 
        p_wishbone_bd_ram_n21467, p_wishbone_bd_ram_n21468, 
        p_wishbone_bd_ram_n21469, p_wishbone_bd_ram_n21470, 
        p_wishbone_bd_ram_n21471, p_wishbone_bd_ram_n21472, 
        p_wishbone_bd_ram_n21473, p_wishbone_bd_ram_n21474, 
        p_wishbone_bd_ram_n21475, p_wishbone_bd_ram_n21476, 
        p_wishbone_bd_ram_n21477, p_wishbone_bd_ram_n21478, 
        p_wishbone_bd_ram_n21479, p_wishbone_bd_ram_n21480, 
        p_wishbone_bd_ram_n21481, p_wishbone_bd_ram_n21482, 
        p_wishbone_bd_ram_n21483, p_wishbone_bd_ram_n21484, 
        p_wishbone_bd_ram_n21485, p_wishbone_bd_ram_n21486, 
        p_wishbone_bd_ram_n21487, p_wishbone_bd_ram_n21488, 
        p_wishbone_bd_ram_n21489, p_wishbone_bd_ram_n21490, 
        p_wishbone_bd_ram_n21491, p_wishbone_bd_ram_n21492, 
        p_wishbone_bd_ram_n21493, p_wishbone_bd_ram_n21494, 
        p_wishbone_bd_ram_n21495, p_wishbone_bd_ram_n21496, 
        p_wishbone_bd_ram_n21497, p_wishbone_bd_ram_n21498, 
        p_wishbone_bd_ram_n21499, p_wishbone_bd_ram_n21500, 
        p_wishbone_bd_ram_n21501, p_wishbone_bd_ram_n21502, 
        p_wishbone_bd_ram_n21503, p_wishbone_bd_ram_n21504, 
        p_wishbone_bd_ram_n21505, p_wishbone_bd_ram_n21506, 
        p_wishbone_bd_ram_n21507, p_wishbone_bd_ram_n21508, 
        p_wishbone_bd_ram_n21509, p_wishbone_bd_ram_n21510, 
        p_wishbone_bd_ram_n21511, p_wishbone_bd_ram_n21512, 
        p_wishbone_bd_ram_n21513, p_wishbone_bd_ram_n21514, 
        p_wishbone_bd_ram_n21515, p_wishbone_bd_ram_n21516, 
        p_wishbone_bd_ram_n21517, p_wishbone_bd_ram_n21518, 
        p_wishbone_bd_ram_n21519, p_wishbone_bd_ram_n21520, 
        p_wishbone_bd_ram_n21521, p_wishbone_bd_ram_n21522, 
        p_wishbone_bd_ram_n21523, p_wishbone_bd_ram_n21524, 
        p_wishbone_bd_ram_n21525, p_wishbone_bd_ram_n21526, 
        p_wishbone_bd_ram_n21527, p_wishbone_bd_ram_n21528, 
        p_wishbone_bd_ram_n21529, p_wishbone_bd_ram_n21530, 
        p_wishbone_bd_ram_n21531, p_wishbone_bd_ram_n21532, 
        p_wishbone_bd_ram_n21533, p_wishbone_bd_ram_n21534, 
        p_wishbone_bd_ram_n21535, p_wishbone_bd_ram_n21536, 
        p_wishbone_bd_ram_n21537, p_wishbone_bd_ram_n21538, 
        p_wishbone_bd_ram_n21539, p_wishbone_bd_ram_n21540, 
        p_wishbone_bd_ram_n21541, p_wishbone_bd_ram_n21542, 
        p_wishbone_bd_ram_n21543, p_wishbone_bd_ram_n21544, 
        p_wishbone_bd_ram_n21545, p_wishbone_bd_ram_n21546, 
        p_wishbone_bd_ram_n21547, p_wishbone_bd_ram_n21548, 
        p_wishbone_bd_ram_n21549, p_wishbone_bd_ram_n21550, 
        p_wishbone_bd_ram_n21551, p_wishbone_bd_ram_n21552, 
        p_wishbone_bd_ram_n21553, p_wishbone_bd_ram_n21554, 
        p_wishbone_bd_ram_n21555, p_wishbone_bd_ram_n21556, 
        p_wishbone_bd_ram_n21557, p_wishbone_bd_ram_n21558, 
        p_wishbone_bd_ram_n21559, p_wishbone_bd_ram_n21560, 
        p_wishbone_bd_ram_n21561, p_wishbone_bd_ram_n21562, 
        p_wishbone_bd_ram_n21563, p_wishbone_bd_ram_n21564, 
        p_wishbone_bd_ram_n21565, p_wishbone_bd_ram_n21566, 
        p_wishbone_bd_ram_n21567, p_wishbone_bd_ram_n21568, 
        p_wishbone_bd_ram_n21569, p_wishbone_bd_ram_n21570, 
        p_wishbone_bd_ram_n21571, p_wishbone_bd_ram_n21572, 
        p_wishbone_bd_ram_n21573, p_wishbone_bd_ram_n21574, 
        p_wishbone_bd_ram_n21575, p_wishbone_bd_ram_n21576, 
        p_wishbone_bd_ram_n21577, p_wishbone_bd_ram_n21578, 
        p_wishbone_bd_ram_n21579, p_wishbone_bd_ram_n21580, 
        p_wishbone_bd_ram_n21581, p_wishbone_bd_ram_n21582, 
        p_wishbone_bd_ram_n21583, p_wishbone_bd_ram_n21584, 
        p_wishbone_bd_ram_n21585, p_wishbone_bd_ram_n21586, 
        p_wishbone_bd_ram_n21587, p_wishbone_bd_ram_n21588, 
        p_wishbone_bd_ram_n21589, p_wishbone_bd_ram_n21590, 
        p_wishbone_bd_ram_n21591, p_wishbone_bd_ram_n21592, 
        p_wishbone_bd_ram_n21593, p_wishbone_bd_ram_n21594, 
        p_wishbone_bd_ram_n21595, p_wishbone_bd_ram_n21596, 
        p_wishbone_bd_ram_n21597, p_wishbone_bd_ram_n21598, 
        p_wishbone_bd_ram_n21599, p_wishbone_bd_ram_n21600, 
        p_wishbone_bd_ram_n21601, p_wishbone_bd_ram_n21602, 
        p_wishbone_bd_ram_n21603, p_wishbone_bd_ram_n21604, 
        p_wishbone_bd_ram_n21605, p_wishbone_bd_ram_n21606, 
        p_wishbone_bd_ram_n21607, p_wishbone_bd_ram_n21608, 
        p_wishbone_bd_ram_n21609, p_wishbone_bd_ram_n21610, 
        p_wishbone_bd_ram_n21611, p_wishbone_bd_ram_n21612, 
        p_wishbone_bd_ram_n21613, p_wishbone_bd_ram_n21614, 
        p_wishbone_bd_ram_n21615, p_wishbone_bd_ram_n21616, 
        p_wishbone_bd_ram_n21617, p_wishbone_bd_ram_n21618, 
        p_wishbone_bd_ram_n21619, p_wishbone_bd_ram_n21620, 
        p_wishbone_bd_ram_n21621, p_wishbone_bd_ram_n21622, 
        p_wishbone_bd_ram_n21623, p_wishbone_bd_ram_n21624, 
        p_wishbone_bd_ram_n21625, p_wishbone_bd_ram_n21626, 
        p_wishbone_bd_ram_n21627, p_wishbone_bd_ram_n21628, 
        p_wishbone_bd_ram_n21629, p_wishbone_bd_ram_n21630, 
        p_wishbone_bd_ram_n21631, p_wishbone_bd_ram_n21632, 
        p_wishbone_bd_ram_n21633, p_wishbone_bd_ram_n21634, 
        p_wishbone_bd_ram_n21635, p_wishbone_bd_ram_n21636, 
        p_wishbone_bd_ram_n21637, p_wishbone_bd_ram_n21638, 
        p_wishbone_bd_ram_n21639, p_wishbone_bd_ram_n21640, 
        p_wishbone_bd_ram_n21641, p_wishbone_bd_ram_n21642, 
        p_wishbone_bd_ram_n21643, p_wishbone_bd_ram_n21644, 
        p_wishbone_bd_ram_n21645, p_wishbone_bd_ram_n21646, 
        p_wishbone_bd_ram_n21647, p_wishbone_bd_ram_n21648, 
        p_wishbone_bd_ram_n21649, p_wishbone_bd_ram_n21650, 
        p_wishbone_bd_ram_n21651, p_wishbone_bd_ram_n21652, 
        p_wishbone_bd_ram_n21653, p_wishbone_bd_ram_n21654, 
        p_wishbone_bd_ram_n21655, p_wishbone_bd_ram_n21656, 
        p_wishbone_bd_ram_n21657, p_wishbone_bd_ram_n21658, 
        p_wishbone_bd_ram_n21659, p_wishbone_bd_ram_n21660, 
        p_wishbone_bd_ram_n21661, p_wishbone_bd_ram_n21662, 
        p_wishbone_bd_ram_n21663, p_wishbone_bd_ram_n21664, 
        p_wishbone_bd_ram_n21665, p_wishbone_bd_ram_n21666, 
        p_wishbone_bd_ram_n21667, p_wishbone_bd_ram_n21668, 
        p_wishbone_bd_ram_n21669, p_wishbone_bd_ram_n21670, 
        p_wishbone_bd_ram_n21671, p_wishbone_bd_ram_n21672, 
        p_wishbone_bd_ram_n21673, p_wishbone_bd_ram_n21674, 
        p_wishbone_bd_ram_n21675, p_wishbone_bd_ram_n21676, 
        p_wishbone_bd_ram_n21677, p_wishbone_bd_ram_n21678, 
        p_wishbone_bd_ram_n21679, p_wishbone_bd_ram_n21680, 
        p_wishbone_bd_ram_n21681, p_wishbone_bd_ram_n21682, 
        p_wishbone_bd_ram_n21683, p_wishbone_bd_ram_n21684, 
        p_wishbone_bd_ram_n21685, p_wishbone_bd_ram_n21686, 
        p_wishbone_bd_ram_n21687, p_wishbone_bd_ram_n21688, 
        p_wishbone_bd_ram_n21689, p_wishbone_bd_ram_n21690, 
        p_wishbone_bd_ram_n21691, p_wishbone_bd_ram_n21692, 
        p_wishbone_bd_ram_n21693, p_wishbone_bd_ram_n21694, 
        p_wishbone_bd_ram_n21695, p_wishbone_bd_ram_n21696, 
        p_wishbone_bd_ram_n21697, p_wishbone_bd_ram_n21698, 
        p_wishbone_bd_ram_n21699, p_wishbone_bd_ram_n21700, 
        p_wishbone_bd_ram_n21701, p_wishbone_bd_ram_n21702, 
        p_wishbone_bd_ram_n21703, p_wishbone_bd_ram_n21704, 
        p_wishbone_bd_ram_n21705, p_wishbone_bd_ram_n21706, 
        p_wishbone_bd_ram_n21707, p_wishbone_bd_ram_n21708, 
        p_wishbone_bd_ram_n21709, p_wishbone_bd_ram_n21710, 
        p_wishbone_bd_ram_n21711, p_wishbone_bd_ram_n21712, 
        p_wishbone_bd_ram_n21713, p_wishbone_bd_ram_n21714, 
        p_wishbone_bd_ram_n21715, p_wishbone_bd_ram_n21716, 
        p_wishbone_bd_ram_n21717, p_wishbone_bd_ram_n21718, 
        p_wishbone_bd_ram_n21719, p_wishbone_bd_ram_n21720, 
        p_wishbone_bd_ram_n21721, p_wishbone_bd_ram_n21722, 
        p_wishbone_bd_ram_n21723, p_wishbone_bd_ram_n21724, 
        p_wishbone_bd_ram_n21725, p_wishbone_bd_ram_n21726, 
        p_wishbone_bd_ram_n21727, p_wishbone_bd_ram_n21728, 
        p_wishbone_bd_ram_n21729, p_wishbone_bd_ram_n21730, 
        p_wishbone_bd_ram_n21731, p_wishbone_bd_ram_n21732, 
        p_wishbone_bd_ram_n21733, p_wishbone_bd_ram_n21734, 
        p_wishbone_bd_ram_n21735, p_wishbone_bd_ram_n21736, 
        p_wishbone_bd_ram_n21737, p_wishbone_bd_ram_n21738, 
        p_wishbone_bd_ram_n21739, p_wishbone_bd_ram_n21740, 
        p_wishbone_bd_ram_n21741, p_wishbone_bd_ram_n21742, 
        p_wishbone_bd_ram_n21743, p_wishbone_bd_ram_n21744, 
        p_wishbone_bd_ram_n21745, p_wishbone_bd_ram_n21746, 
        p_wishbone_bd_ram_n21747, p_wishbone_bd_ram_n21748, 
        p_wishbone_bd_ram_n21749, p_wishbone_bd_ram_n21750, 
        p_wishbone_bd_ram_n21751, p_wishbone_bd_ram_n21752, 
        p_wishbone_bd_ram_n21753, p_wishbone_bd_ram_n21754, 
        p_wishbone_bd_ram_n21755, p_wishbone_bd_ram_n21756, 
        p_wishbone_bd_ram_n21757, p_wishbone_bd_ram_n21758, 
        p_wishbone_bd_ram_n21759, p_wishbone_bd_ram_n21760, 
        p_wishbone_bd_ram_n21761, p_wishbone_bd_ram_n21762, 
        p_wishbone_bd_ram_n21763, p_wishbone_bd_ram_n21764, 
        p_wishbone_bd_ram_n21765, p_wishbone_bd_ram_n21766, 
        p_wishbone_bd_ram_n21767, p_wishbone_bd_ram_n21768, 
        p_wishbone_bd_ram_n21769, p_wishbone_bd_ram_n21770, 
        p_wishbone_bd_ram_n21771, p_wishbone_bd_ram_n21772, 
        p_wishbone_bd_ram_n21773, p_wishbone_bd_ram_n21774, 
        p_wishbone_bd_ram_n21775, p_wishbone_bd_ram_n21776, 
        p_wishbone_bd_ram_n21777, p_wishbone_bd_ram_n21778, 
        p_wishbone_bd_ram_n21779, p_wishbone_bd_ram_n21780, 
        p_wishbone_bd_ram_n21781, p_wishbone_bd_ram_n21782, 
        p_wishbone_bd_ram_n21783, p_wishbone_bd_ram_n21784, 
        p_wishbone_bd_ram_n21785, p_wishbone_bd_ram_n21786, 
        p_wishbone_bd_ram_n21787, p_wishbone_bd_ram_n21788, 
        p_wishbone_bd_ram_n21789, p_wishbone_bd_ram_n21790, 
        p_wishbone_bd_ram_n21791, p_wishbone_bd_ram_n21792, 
        p_wishbone_bd_ram_n21793, p_wishbone_bd_ram_n21794, 
        p_wishbone_bd_ram_n21795, p_wishbone_bd_ram_n21796, 
        p_wishbone_bd_ram_n21797, p_wishbone_bd_ram_n21798, 
        p_wishbone_bd_ram_n21799, p_wishbone_bd_ram_n21800, 
        p_wishbone_bd_ram_n21801, p_wishbone_bd_ram_n21802, 
        p_wishbone_bd_ram_n21803, p_wishbone_bd_ram_n21804, 
        p_wishbone_bd_ram_n21805, p_wishbone_bd_ram_n21806, 
        p_wishbone_bd_ram_n21807, p_wishbone_bd_ram_n21808, 
        p_wishbone_bd_ram_n21809, p_wishbone_bd_ram_n21810, 
        p_wishbone_bd_ram_n21811, p_wishbone_bd_ram_n21812, 
        p_wishbone_bd_ram_n21813, p_wishbone_bd_ram_n21814, 
        p_wishbone_bd_ram_n21815, p_wishbone_bd_ram_n21816, 
        p_wishbone_bd_ram_n21817, p_wishbone_bd_ram_n21818, 
        p_wishbone_bd_ram_n21819, p_wishbone_bd_ram_n21820, 
        p_wishbone_bd_ram_n21821, p_wishbone_bd_ram_n21822, 
        p_wishbone_bd_ram_n21823, p_wishbone_bd_ram_n21824, 
        p_wishbone_bd_ram_n21825, p_wishbone_bd_ram_n21826, 
        p_wishbone_bd_ram_n21827, p_wishbone_bd_ram_n21828, 
        p_wishbone_bd_ram_n21829, p_wishbone_bd_ram_n21830, 
        p_wishbone_bd_ram_n21831, p_wishbone_bd_ram_n21832, 
        p_wishbone_bd_ram_n21833, p_wishbone_bd_ram_n21834, 
        p_wishbone_bd_ram_n21835, p_wishbone_bd_ram_n21836, 
        p_wishbone_bd_ram_n21837, p_wishbone_bd_ram_n21838, 
        p_wishbone_bd_ram_n21839, p_wishbone_bd_ram_n21840, 
        p_wishbone_bd_ram_n21841, p_wishbone_bd_ram_n21842, 
        p_wishbone_bd_ram_n21843, p_wishbone_bd_ram_n21844, 
        p_wishbone_bd_ram_n21845, p_wishbone_bd_ram_n21846, 
        p_wishbone_bd_ram_n21847, p_wishbone_bd_ram_n21848, 
        p_wishbone_bd_ram_n21849, p_wishbone_bd_ram_n21850, 
        p_wishbone_bd_ram_n21851, p_wishbone_bd_ram_n21852, 
        p_wishbone_bd_ram_n21853, p_wishbone_bd_ram_n21854, 
        p_wishbone_bd_ram_n21855, p_wishbone_bd_ram_n21856, 
        p_wishbone_bd_ram_n21857, p_wishbone_bd_ram_n21858, 
        p_wishbone_bd_ram_n21859, p_wishbone_bd_ram_n21860, 
        p_wishbone_bd_ram_n21861, p_wishbone_bd_ram_n21862, 
        p_wishbone_bd_ram_n21863, p_wishbone_bd_ram_n21864, 
        p_wishbone_bd_ram_n21865, p_wishbone_bd_ram_n21866, 
        p_wishbone_bd_ram_n21867, p_wishbone_bd_ram_n21868, 
        p_wishbone_bd_ram_n21869, p_wishbone_bd_ram_n21870, 
        p_wishbone_bd_ram_n21871, p_wishbone_bd_ram_n21872, 
        p_wishbone_bd_ram_n21873, p_wishbone_bd_ram_n21874, 
        p_wishbone_bd_ram_n21875, p_wishbone_bd_ram_n21876, 
        p_wishbone_bd_ram_n21877, p_wishbone_bd_ram_n21878, 
        p_wishbone_bd_ram_n21879, p_wishbone_bd_ram_n21880, 
        p_wishbone_bd_ram_n21881, p_wishbone_bd_ram_n21882, 
        p_wishbone_bd_ram_n21883, p_wishbone_bd_ram_n21884, 
        p_wishbone_bd_ram_n21885, p_wishbone_bd_ram_n21886, 
        p_wishbone_bd_ram_n21887, p_wishbone_bd_ram_n21888, 
        p_wishbone_bd_ram_n21889, p_wishbone_bd_ram_n21890, 
        p_wishbone_bd_ram_n21891, p_wishbone_bd_ram_n21892, 
        p_wishbone_bd_ram_n21893, p_wishbone_bd_ram_n21894, 
        p_wishbone_bd_ram_n21895, p_wishbone_bd_ram_n21896, 
        p_wishbone_bd_ram_n21897, p_wishbone_bd_ram_n21898, 
        p_wishbone_bd_ram_n21899, p_wishbone_bd_ram_n21900, 
        p_wishbone_bd_ram_n21901, p_wishbone_bd_ram_n21902, 
        p_wishbone_bd_ram_n21903, p_wishbone_bd_ram_n21904, 
        p_wishbone_bd_ram_n21905, p_wishbone_bd_ram_n21906, 
        p_wishbone_bd_ram_n21907, p_wishbone_bd_ram_n21908, 
        p_wishbone_bd_ram_n21909, p_wishbone_bd_ram_n21910, 
        p_wishbone_bd_ram_n21911, p_wishbone_bd_ram_n21912, 
        p_wishbone_bd_ram_n21913, p_wishbone_bd_ram_n21914, 
        p_wishbone_bd_ram_n21915, p_wishbone_bd_ram_n21916, 
        p_wishbone_bd_ram_n21917, p_wishbone_bd_ram_n21918, 
        p_wishbone_bd_ram_n21919, p_wishbone_bd_ram_n21920, 
        p_wishbone_bd_ram_n21921, p_wishbone_bd_ram_n21922, 
        p_wishbone_bd_ram_n21923, p_wishbone_bd_ram_n21924, 
        p_wishbone_bd_ram_n21925, p_wishbone_bd_ram_n21926, 
        p_wishbone_bd_ram_n21927, p_wishbone_bd_ram_n21928, 
        p_wishbone_bd_ram_n21929, p_wishbone_bd_ram_n21930, 
        p_wishbone_bd_ram_n21931, p_wishbone_bd_ram_n21932, 
        p_wishbone_bd_ram_n21933, p_wishbone_bd_ram_n21934, 
        p_wishbone_bd_ram_n21935, p_wishbone_bd_ram_n21936, 
        p_wishbone_bd_ram_n21937, p_wishbone_bd_ram_n21938, 
        p_wishbone_bd_ram_n21939, p_wishbone_bd_ram_n21940, 
        p_wishbone_bd_ram_n21941, p_wishbone_bd_ram_n21942, 
        p_wishbone_bd_ram_n21943, p_wishbone_bd_ram_n21944, 
        p_wishbone_bd_ram_n21945, p_wishbone_bd_ram_n21946, 
        p_wishbone_bd_ram_n21947, p_wishbone_bd_ram_n21948, 
        p_wishbone_bd_ram_n21949, p_wishbone_bd_ram_n21950, 
        p_wishbone_bd_ram_n21951, p_wishbone_bd_ram_n21952, 
        p_wishbone_bd_ram_n21953, p_wishbone_bd_ram_n21954, 
        p_wishbone_bd_ram_n21955, p_wishbone_bd_ram_n21956, 
        p_wishbone_bd_ram_n21957, p_wishbone_bd_ram_n21958, 
        p_wishbone_bd_ram_n21959, p_wishbone_bd_ram_n21960, 
        p_wishbone_bd_ram_n21961, p_wishbone_bd_ram_n21962, 
        p_wishbone_bd_ram_n21963, p_wishbone_bd_ram_n21964, 
        p_wishbone_bd_ram_n21965, p_wishbone_bd_ram_n21966, 
        p_wishbone_bd_ram_n21967, p_wishbone_bd_ram_n21968, 
        p_wishbone_bd_ram_n21969, p_wishbone_bd_ram_n21970, 
        p_wishbone_bd_ram_n21971, p_wishbone_bd_ram_n21972, 
        p_wishbone_bd_ram_n21973, p_wishbone_bd_ram_n21974, 
        p_wishbone_bd_ram_n21975, p_wishbone_bd_ram_n21976, 
        p_wishbone_bd_ram_n21977, p_wishbone_bd_ram_n21978, 
        p_wishbone_bd_ram_n21979, p_wishbone_bd_ram_n21980, 
        p_wishbone_bd_ram_n21981, p_wishbone_bd_ram_n21982, 
        p_wishbone_bd_ram_n21983, p_wishbone_bd_ram_n21984, 
        p_wishbone_bd_ram_n21985, p_wishbone_bd_ram_n21986, 
        p_wishbone_bd_ram_n21987, p_wishbone_bd_ram_n21988, 
        p_wishbone_bd_ram_n21989, p_wishbone_bd_ram_n21990, 
        p_wishbone_bd_ram_n21991, p_wishbone_bd_ram_n21992, 
        p_wishbone_bd_ram_n21993, p_wishbone_bd_ram_n21994, 
        p_wishbone_bd_ram_n21995, p_wishbone_bd_ram_n21996, 
        p_wishbone_bd_ram_n21997, p_wishbone_bd_ram_n21998, 
        p_wishbone_bd_ram_n21999, p_wishbone_bd_ram_n22000, 
        p_wishbone_bd_ram_n22001, p_wishbone_bd_ram_n22002, 
        p_wishbone_bd_ram_n22003, p_wishbone_bd_ram_n22004, 
        p_wishbone_bd_ram_n22005, p_wishbone_bd_ram_n22006, 
        p_wishbone_bd_ram_n22007, p_wishbone_bd_ram_n22008, 
        p_wishbone_bd_ram_n22009, p_wishbone_bd_ram_n22010, 
        p_wishbone_bd_ram_n22011, p_wishbone_bd_ram_n22012, 
        p_wishbone_bd_ram_n22013, p_wishbone_bd_ram_n22014, 
        p_wishbone_bd_ram_n22015, p_wishbone_bd_ram_n22016, 
        p_wishbone_bd_ram_n22017, p_wishbone_bd_ram_n22018, 
        p_wishbone_bd_ram_n22019, p_wishbone_bd_ram_n22020, 
        p_wishbone_bd_ram_n22021, p_wishbone_bd_ram_n22022, 
        p_wishbone_bd_ram_n22023, p_wishbone_bd_ram_n22024, 
        p_wishbone_bd_ram_n22025, p_wishbone_bd_ram_n22026, 
        p_wishbone_bd_ram_n22027, p_wishbone_bd_ram_n22028, 
        p_wishbone_bd_ram_n22029, p_wishbone_bd_ram_n22030, 
        p_wishbone_bd_ram_n22031, p_wishbone_bd_ram_n22032, 
        p_wishbone_bd_ram_n22033, p_wishbone_bd_ram_n22034, 
        p_wishbone_bd_ram_n22035, p_wishbone_bd_ram_n22036, 
        p_wishbone_bd_ram_n22037, p_wishbone_bd_ram_n22038, 
        p_wishbone_bd_ram_n22039, p_wishbone_bd_ram_n22040, 
        p_wishbone_bd_ram_n22041, p_wishbone_bd_ram_n22042, 
        p_wishbone_bd_ram_n22043, p_wishbone_bd_ram_n22044, 
        p_wishbone_bd_ram_n22045, p_wishbone_bd_ram_n22046, 
        p_wishbone_bd_ram_n22047, p_wishbone_bd_ram_n22048, 
        p_wishbone_bd_ram_n22049, p_wishbone_bd_ram_n22050, 
        p_wishbone_bd_ram_n22051, p_wishbone_bd_ram_n22052, 
        p_wishbone_bd_ram_n22053, p_wishbone_bd_ram_n22054, 
        p_wishbone_bd_ram_n22055, p_wishbone_bd_ram_n22056, 
        p_wishbone_bd_ram_n22057, p_wishbone_bd_ram_n22058, 
        p_wishbone_bd_ram_n22059, p_wishbone_bd_ram_n22060, 
        p_wishbone_bd_ram_n22061, p_wishbone_bd_ram_n22062, 
        p_wishbone_bd_ram_n22063, p_wishbone_bd_ram_n22064, 
        p_wishbone_bd_ram_n22065, p_wishbone_bd_ram_n22066, 
        p_wishbone_bd_ram_n22067, p_wishbone_bd_ram_n22068, 
        p_wishbone_bd_ram_n22069, p_wishbone_bd_ram_n22070, 
        p_wishbone_bd_ram_n22071, p_wishbone_bd_ram_n22072, 
        p_wishbone_bd_ram_n22073, p_wishbone_bd_ram_n22074, 
        p_wishbone_bd_ram_n22075, p_wishbone_bd_ram_n22076, 
        p_wishbone_bd_ram_n22077, p_wishbone_bd_ram_n22078, 
        p_wishbone_bd_ram_n22079, p_wishbone_bd_ram_n22080, 
        p_wishbone_bd_ram_n22081, p_wishbone_bd_ram_n22082, 
        p_wishbone_bd_ram_n22083, p_wishbone_bd_ram_n22084, 
        p_wishbone_bd_ram_n22085, p_wishbone_bd_ram_n22086, 
        p_wishbone_bd_ram_n22087, p_wishbone_bd_ram_n22088, 
        p_wishbone_bd_ram_n22089, p_wishbone_bd_ram_n22090, 
        p_wishbone_bd_ram_n22091, p_wishbone_bd_ram_n22092, 
        p_wishbone_bd_ram_n22093, p_wishbone_bd_ram_n22094, 
        p_wishbone_bd_ram_n22095, p_wishbone_bd_ram_n22096, 
        p_wishbone_bd_ram_n22097, p_wishbone_bd_ram_n22098, 
        p_wishbone_bd_ram_n22099, p_wishbone_bd_ram_n22100, 
        p_wishbone_bd_ram_n22101, p_wishbone_bd_ram_n22102, 
        p_wishbone_bd_ram_n22103, p_wishbone_bd_ram_n22104, 
        p_wishbone_bd_ram_n22105, p_wishbone_bd_ram_n22106, 
        p_wishbone_bd_ram_n22107, p_wishbone_bd_ram_n22108, 
        p_wishbone_bd_ram_n22109, p_wishbone_bd_ram_n22110, 
        p_wishbone_bd_ram_n22111, p_wishbone_bd_ram_n22112, 
        p_wishbone_bd_ram_n22113, p_wishbone_bd_ram_n22114, 
        p_wishbone_bd_ram_n22115, p_wishbone_bd_ram_n22116, 
        p_wishbone_bd_ram_n22117, p_wishbone_bd_ram_n22118, 
        p_wishbone_bd_ram_n22119, p_wishbone_bd_ram_n22120, 
        p_wishbone_bd_ram_n22121, p_wishbone_bd_ram_n22122, 
        p_wishbone_bd_ram_n22123, p_wishbone_bd_ram_n22124, 
        p_wishbone_bd_ram_n22125, p_wishbone_bd_ram_n22126, 
        p_wishbone_bd_ram_n22127, p_wishbone_bd_ram_n22128, 
        p_wishbone_bd_ram_n22129, p_wishbone_bd_ram_n22130, 
        p_wishbone_bd_ram_n22131, p_wishbone_bd_ram_n22132, 
        p_wishbone_bd_ram_n22133, p_wishbone_bd_ram_n22134, 
        p_wishbone_bd_ram_n22135, p_wishbone_bd_ram_n22136, 
        p_wishbone_bd_ram_n22137, p_wishbone_bd_ram_n22138, 
        p_wishbone_bd_ram_n22139, p_wishbone_bd_ram_n22140, 
        p_wishbone_bd_ram_n22141, p_wishbone_bd_ram_n22142, 
        p_wishbone_bd_ram_n22143, p_wishbone_bd_ram_n22144, 
        p_wishbone_bd_ram_n22145, p_wishbone_bd_ram_n22146, 
        p_wishbone_bd_ram_n22147, p_wishbone_bd_ram_n22148, 
        p_wishbone_bd_ram_n22149, p_wishbone_bd_ram_n22150, 
        p_wishbone_bd_ram_n22151, p_wishbone_bd_ram_n22152, 
        p_wishbone_bd_ram_n22153, p_wishbone_bd_ram_n22154, 
        p_wishbone_bd_ram_n22155, p_wishbone_bd_ram_n22156, 
        p_wishbone_bd_ram_n22157, p_wishbone_bd_ram_n22158, 
        p_wishbone_bd_ram_n22159, p_wishbone_bd_ram_n22160, 
        p_wishbone_bd_ram_n22161, p_wishbone_bd_ram_n22162, 
        p_wishbone_bd_ram_n22163, p_wishbone_bd_ram_n22164, 
        p_wishbone_bd_ram_n22165, p_wishbone_bd_ram_n22166, 
        p_wishbone_bd_ram_n22167, p_wishbone_bd_ram_n22168, 
        p_wishbone_bd_ram_n22169, p_wishbone_bd_ram_n22170, 
        p_wishbone_bd_ram_n22171, p_wishbone_bd_ram_n22172, 
        p_wishbone_bd_ram_n22173, p_wishbone_bd_ram_n22174, 
        p_wishbone_bd_ram_n22175, p_wishbone_bd_ram_n22176, 
        p_wishbone_bd_ram_n22177, p_wishbone_bd_ram_n22178, 
        p_wishbone_bd_ram_n22179, p_wishbone_bd_ram_n22180, 
        p_wishbone_bd_ram_n22181, p_wishbone_bd_ram_n22182, 
        p_wishbone_bd_ram_n22183, p_wishbone_bd_ram_n22184, 
        p_wishbone_bd_ram_n22185, p_wishbone_bd_ram_n22186, 
        p_wishbone_bd_ram_n22187, p_wishbone_bd_ram_n22188, 
        p_wishbone_bd_ram_n22189, p_wishbone_bd_ram_n22190, 
        p_wishbone_bd_ram_n22191, p_wishbone_bd_ram_n22192, 
        p_wishbone_bd_ram_n22193, p_wishbone_bd_ram_n22194, 
        p_wishbone_bd_ram_n22195, p_wishbone_bd_ram_n22196, 
        p_wishbone_bd_ram_n22197, p_wishbone_bd_ram_n22198, 
        p_wishbone_bd_ram_n22199, p_wishbone_bd_ram_n22200, 
        p_wishbone_bd_ram_n22201, p_wishbone_bd_ram_n22202, 
        p_wishbone_bd_ram_n22203, p_wishbone_bd_ram_n22204, 
        p_wishbone_bd_ram_n22205, p_wishbone_bd_ram_n22206, 
        p_wishbone_bd_ram_n22207, p_wishbone_bd_ram_n22208, 
        p_wishbone_bd_ram_n22209, p_wishbone_bd_ram_n22210, 
        p_wishbone_bd_ram_n22211, p_wishbone_bd_ram_n22212, 
        p_wishbone_bd_ram_n22213, p_wishbone_bd_ram_n22214, 
        p_wishbone_bd_ram_n22215, p_wishbone_bd_ram_n22216, 
        p_wishbone_bd_ram_n22217, p_wishbone_bd_ram_n22218, 
        p_wishbone_bd_ram_n22219, p_wishbone_bd_ram_n22220, 
        p_wishbone_bd_ram_n22221, p_wishbone_bd_ram_n22222, 
        p_wishbone_bd_ram_n22223, p_wishbone_bd_ram_n22224, 
        p_wishbone_bd_ram_n22225, p_wishbone_bd_ram_n22226, 
        p_wishbone_bd_ram_n22227, p_wishbone_bd_ram_n22228, 
        p_wishbone_bd_ram_n22229, p_wishbone_bd_ram_n22230, 
        p_wishbone_bd_ram_n22231, p_wishbone_bd_ram_n22232, 
        p_wishbone_bd_ram_n22233, p_wishbone_bd_ram_n22234, 
        p_wishbone_bd_ram_n22235, p_wishbone_bd_ram_n22236, 
        p_wishbone_bd_ram_n22237, p_wishbone_bd_ram_n22238, 
        p_wishbone_bd_ram_n22239, p_wishbone_bd_ram_n22240, 
        p_wishbone_bd_ram_n22241, p_wishbone_bd_ram_n22242, 
        p_wishbone_bd_ram_n22243, p_wishbone_bd_ram_n22244, 
        p_wishbone_bd_ram_n22245, p_wishbone_bd_ram_n22246, 
        p_wishbone_bd_ram_n22247, p_wishbone_bd_ram_n22248, 
        p_wishbone_bd_ram_n22249, p_wishbone_bd_ram_n22250, 
        p_wishbone_bd_ram_n22251, p_wishbone_bd_ram_n22252, 
        p_wishbone_bd_ram_n22253, p_wishbone_bd_ram_n22254, 
        p_wishbone_bd_ram_n22255, p_wishbone_bd_ram_n22256, 
        p_wishbone_bd_ram_n22257, p_wishbone_bd_ram_n22258, 
        p_wishbone_bd_ram_n22259, p_wishbone_bd_ram_n22260, 
        p_wishbone_bd_ram_n22261, p_wishbone_bd_ram_n22262, 
        p_wishbone_bd_ram_n22263, p_wishbone_bd_ram_n22264, 
        p_wishbone_bd_ram_n22265, p_wishbone_bd_ram_n22266, 
        p_wishbone_bd_ram_n22267, p_wishbone_bd_ram_n22268, 
        p_wishbone_bd_ram_n22269, p_wishbone_bd_ram_n22270, 
        p_wishbone_bd_ram_n22271, p_wishbone_bd_ram_n22272, 
        p_wishbone_bd_ram_n22273, p_wishbone_bd_ram_n22274, 
        p_wishbone_bd_ram_n22275, p_wishbone_bd_ram_n22276, 
        p_wishbone_bd_ram_n22277, p_wishbone_bd_ram_n22278, 
        p_wishbone_bd_ram_n22279, p_wishbone_bd_ram_n22280, 
        p_wishbone_bd_ram_n22281, p_wishbone_bd_ram_n22282, 
        p_wishbone_bd_ram_n22283, p_wishbone_bd_ram_n22284, 
        p_wishbone_bd_ram_n22285, p_wishbone_bd_ram_n22286, 
        p_wishbone_bd_ram_n22287, p_wishbone_bd_ram_n22288, 
        p_wishbone_bd_ram_n22289, p_wishbone_bd_ram_n22290, 
        p_wishbone_bd_ram_n22291, p_wishbone_bd_ram_n22292, 
        p_wishbone_bd_ram_n22293, p_wishbone_bd_ram_n22294, 
        p_wishbone_bd_ram_n22295, p_wishbone_bd_ram_n22296, 
        p_wishbone_bd_ram_n22297, p_wishbone_bd_ram_n22298, 
        p_wishbone_bd_ram_n22299, p_wishbone_bd_ram_n22300, 
        p_wishbone_bd_ram_n22301, p_wishbone_bd_ram_n22302, 
        p_wishbone_bd_ram_n22303, p_wishbone_bd_ram_n22304, 
        p_wishbone_bd_ram_n22305, p_wishbone_bd_ram_n22306, 
        p_wishbone_bd_ram_n22307, p_wishbone_bd_ram_n22308, 
        p_wishbone_bd_ram_n22309, p_wishbone_bd_ram_n22310, 
        p_wishbone_bd_ram_n22311, p_wishbone_bd_ram_n22312, 
        p_wishbone_bd_ram_n22313, p_wishbone_bd_ram_n22314, 
        p_wishbone_bd_ram_n22315, p_wishbone_bd_ram_n22316, 
        p_wishbone_bd_ram_n22317, p_wishbone_bd_ram_n22318, 
        p_wishbone_bd_ram_n22319, p_wishbone_bd_ram_n22320, 
        p_wishbone_bd_ram_n22321, p_wishbone_bd_ram_n22322, 
        p_wishbone_bd_ram_n22323, p_wishbone_bd_ram_n22324, 
        p_wishbone_bd_ram_n22325, p_wishbone_bd_ram_n22326, 
        p_wishbone_bd_ram_n22327, p_wishbone_bd_ram_n22328, 
        p_wishbone_bd_ram_n22329, p_wishbone_bd_ram_n22330, 
        p_wishbone_bd_ram_n22331, p_wishbone_bd_ram_n22332, 
        p_wishbone_bd_ram_n22333, p_wishbone_bd_ram_n22334, 
        p_wishbone_bd_ram_n22335, p_wishbone_bd_ram_n22336, 
        p_wishbone_bd_ram_n22337, p_wishbone_bd_ram_n22338, 
        p_wishbone_bd_ram_n22339, p_wishbone_bd_ram_n22340, 
        p_wishbone_bd_ram_n22341, p_wishbone_bd_ram_n22342, 
        p_wishbone_bd_ram_n22343, p_wishbone_bd_ram_n22344, 
        p_wishbone_bd_ram_n22345, p_wishbone_bd_ram_n22346, 
        p_wishbone_bd_ram_n22347, p_wishbone_bd_ram_n22348, 
        p_wishbone_bd_ram_n22349, p_wishbone_bd_ram_n22350, 
        p_wishbone_bd_ram_n22351, p_wishbone_bd_ram_n22352, 
        p_wishbone_bd_ram_n22353, p_wishbone_bd_ram_n22354, 
        p_wishbone_bd_ram_n22355, p_wishbone_bd_ram_n22356, 
        p_wishbone_bd_ram_n22357, p_wishbone_bd_ram_n22358, 
        p_wishbone_bd_ram_n22359, p_wishbone_bd_ram_n22360, 
        p_wishbone_bd_ram_n22361, p_wishbone_bd_ram_n22362, 
        p_wishbone_bd_ram_n22363, p_wishbone_bd_ram_n22364, 
        p_wishbone_bd_ram_n22365, p_wishbone_bd_ram_n22366, 
        p_wishbone_bd_ram_n22367, p_wishbone_bd_ram_n22368, 
        p_wishbone_bd_ram_n22369, p_wishbone_bd_ram_n22370, 
        p_wishbone_bd_ram_n22371, p_wishbone_bd_ram_n22372, 
        p_wishbone_bd_ram_n22373, p_wishbone_bd_ram_n22374, 
        p_wishbone_bd_ram_n22375, p_wishbone_bd_ram_n22376, 
        p_wishbone_bd_ram_n22377, p_wishbone_bd_ram_n22378, 
        p_wishbone_bd_ram_n22379, p_wishbone_bd_ram_n22380, 
        p_wishbone_bd_ram_n22381, p_wishbone_bd_ram_n22382, 
        p_wishbone_bd_ram_n22383, p_wishbone_bd_ram_n22384, 
        p_wishbone_bd_ram_n22385, p_wishbone_bd_ram_n22386, 
        p_wishbone_bd_ram_n22387, p_wishbone_bd_ram_n22388, 
        p_wishbone_bd_ram_n22389, p_wishbone_bd_ram_n22390, 
        p_wishbone_bd_ram_n22391, p_wishbone_bd_ram_n22392, 
        p_wishbone_bd_ram_n22393, p_wishbone_bd_ram_n22394, 
        p_wishbone_bd_ram_n22395, p_wishbone_bd_ram_n22396, 
        p_wishbone_bd_ram_n22397, p_wishbone_bd_ram_n22398, 
        p_wishbone_bd_ram_n22399, p_wishbone_bd_ram_n22400, 
        p_wishbone_bd_ram_n22401, p_wishbone_bd_ram_n22402, 
        p_wishbone_bd_ram_n22403, p_wishbone_bd_ram_n22404, 
        p_wishbone_bd_ram_n22405, p_wishbone_bd_ram_n22406, 
        p_wishbone_bd_ram_n22407, p_wishbone_bd_ram_n22408, 
        p_wishbone_bd_ram_n22409, p_wishbone_bd_ram_n22410, 
        p_wishbone_bd_ram_n22411, p_wishbone_bd_ram_n22412, 
        p_wishbone_bd_ram_n22413, p_wishbone_bd_ram_n22414, 
        p_wishbone_bd_ram_n22415, p_wishbone_bd_ram_n22416, 
        p_wishbone_bd_ram_n22417, p_wishbone_bd_ram_n22418, 
        p_wishbone_bd_ram_n22419, p_wishbone_bd_ram_n22420, 
        p_wishbone_bd_ram_n22421, p_wishbone_bd_ram_n22422, 
        p_wishbone_bd_ram_n22423, p_wishbone_bd_ram_n22424, 
        p_wishbone_bd_ram_n22425, p_wishbone_bd_ram_n22426, 
        p_wishbone_bd_ram_n22427, p_wishbone_bd_ram_n22428, 
        p_wishbone_bd_ram_n22429, p_wishbone_bd_ram_n22430, 
        p_wishbone_bd_ram_n22431, p_wishbone_bd_ram_n22432, 
        p_wishbone_bd_ram_n22433, p_wishbone_bd_ram_n22434, 
        p_wishbone_bd_ram_n22435, p_wishbone_bd_ram_n22436, 
        p_wishbone_bd_ram_n22437, p_wishbone_bd_ram_n22438, 
        p_wishbone_bd_ram_n22439, p_wishbone_bd_ram_n22440, 
        p_wishbone_bd_ram_n22441, p_wishbone_bd_ram_n22442, 
        p_wishbone_bd_ram_n22443, p_wishbone_bd_ram_n22444, 
        p_wishbone_bd_ram_n22445, p_wishbone_bd_ram_n22446, 
        p_wishbone_bd_ram_n22447, p_wishbone_bd_ram_n22448, 
        p_wishbone_bd_ram_n22449, p_wishbone_bd_ram_n22450, 
        p_wishbone_bd_ram_n22451, p_wishbone_bd_ram_n22452, 
        p_wishbone_bd_ram_n22453, p_wishbone_bd_ram_n22454, 
        p_wishbone_bd_ram_n22455, p_wishbone_bd_ram_n22456, 
        p_wishbone_bd_ram_n22457, p_wishbone_bd_ram_n22458, 
        p_wishbone_bd_ram_n22459, p_wishbone_bd_ram_n22460, 
        p_wishbone_bd_ram_n22461, p_wishbone_bd_ram_n22462, 
        p_wishbone_bd_ram_n22463, p_wishbone_bd_ram_n22464, 
        p_wishbone_bd_ram_n22465, p_wishbone_bd_ram_n22466, 
        p_wishbone_bd_ram_n22467, p_wishbone_bd_ram_n22468, 
        p_wishbone_bd_ram_n22469, p_wishbone_bd_ram_n22470, 
        p_wishbone_bd_ram_n22471, p_wishbone_bd_ram_n22472, 
        p_wishbone_bd_ram_n22473, p_wishbone_bd_ram_n22474, 
        p_wishbone_bd_ram_n22475, p_wishbone_bd_ram_n22476, 
        p_wishbone_bd_ram_n22477, p_wishbone_bd_ram_n22478, 
        p_wishbone_bd_ram_n22479, p_wishbone_bd_ram_n22480, 
        p_wishbone_bd_ram_n22481, p_wishbone_bd_ram_n22482, 
        p_wishbone_bd_ram_n22483, p_wishbone_bd_ram_n22484, 
        p_wishbone_bd_ram_n22485, p_wishbone_bd_ram_n22486, 
        p_wishbone_bd_ram_n22487, p_wishbone_bd_ram_n22488, 
        p_wishbone_bd_ram_n22489, p_wishbone_bd_ram_n22490, 
        p_wishbone_bd_ram_n22491, p_wishbone_bd_ram_n22492, 
        p_wishbone_bd_ram_n22493, p_wishbone_bd_ram_n22494, 
        p_wishbone_bd_ram_n22495, p_wishbone_bd_ram_n22496, 
        p_wishbone_bd_ram_n22497, p_wishbone_bd_ram_n22498, 
        p_wishbone_bd_ram_n22499, p_wishbone_bd_ram_n22500, 
        p_wishbone_bd_ram_n22501, p_wishbone_bd_ram_n22502, 
        p_wishbone_bd_ram_n22503, p_wishbone_bd_ram_n22504, 
        p_wishbone_bd_ram_n22505, p_wishbone_bd_ram_n22506, 
        p_wishbone_bd_ram_n22507, p_wishbone_bd_ram_n22508, 
        p_wishbone_bd_ram_n22509, p_wishbone_bd_ram_n22510, 
        p_wishbone_bd_ram_n22511, p_wishbone_bd_ram_n22512, 
        p_wishbone_bd_ram_n22513, p_wishbone_bd_ram_n22514, 
        p_wishbone_bd_ram_n22515, p_wishbone_bd_ram_n22516, 
        p_wishbone_bd_ram_n22517, p_wishbone_bd_ram_n22518, 
        p_wishbone_bd_ram_n22519, p_wishbone_bd_ram_n22520, 
        p_wishbone_bd_ram_n22521, p_wishbone_bd_ram_n22522, 
        p_wishbone_bd_ram_n22523, p_wishbone_bd_ram_n22524, 
        p_wishbone_bd_ram_n22525, p_wishbone_bd_ram_n22526, 
        p_wishbone_bd_ram_n22527, p_wishbone_bd_ram_n22528, 
        p_wishbone_bd_ram_n22529, p_wishbone_bd_ram_n22530, 
        p_wishbone_bd_ram_n22531, p_wishbone_bd_ram_n22532, 
        p_wishbone_bd_ram_n22533, p_wishbone_bd_ram_n22534, 
        p_wishbone_bd_ram_n22535, p_wishbone_bd_ram_n22536, 
        p_wishbone_bd_ram_n22537, p_wishbone_bd_ram_n22538, 
        p_wishbone_bd_ram_n22539, p_wishbone_bd_ram_n22540, 
        p_wishbone_bd_ram_n22541, p_wishbone_bd_ram_n22542, 
        p_wishbone_bd_ram_n22543, p_wishbone_bd_ram_n22544, 
        p_wishbone_bd_ram_n22545, p_wishbone_bd_ram_n22546, 
        p_wishbone_bd_ram_n22547, p_wishbone_bd_ram_n22548, 
        p_wishbone_bd_ram_n22549, p_wishbone_bd_ram_n22550, 
        p_wishbone_bd_ram_n22551, p_wishbone_bd_ram_n22552, 
        p_wishbone_bd_ram_n22553, p_wishbone_bd_ram_n22554, 
        p_wishbone_bd_ram_n22555, p_wishbone_bd_ram_n22556, 
        p_wishbone_bd_ram_n22557, p_wishbone_bd_ram_n22558, 
        p_wishbone_bd_ram_n22559, p_wishbone_bd_ram_n22560, 
        p_wishbone_bd_ram_n22561, p_wishbone_bd_ram_n22562, 
        p_wishbone_bd_ram_n22563, p_wishbone_bd_ram_n22564, 
        p_wishbone_bd_ram_n22565, p_wishbone_bd_ram_n22566, 
        p_wishbone_bd_ram_n22567, p_wishbone_bd_ram_n22568, 
        p_wishbone_bd_ram_n22569, p_wishbone_bd_ram_n22570, 
        p_wishbone_bd_ram_n22571, p_wishbone_bd_ram_n22572, 
        p_wishbone_bd_ram_n22573, p_wishbone_bd_ram_n22574, 
        p_wishbone_bd_ram_n22575, p_wishbone_bd_ram_n22576, 
        p_wishbone_bd_ram_n22577, p_wishbone_bd_ram_n22578, 
        p_wishbone_bd_ram_n22579, p_wishbone_bd_ram_n22580, 
        p_wishbone_bd_ram_n22581, p_wishbone_bd_ram_n22582, 
        p_wishbone_bd_ram_n22583, p_wishbone_bd_ram_n22584, 
        p_wishbone_bd_ram_n22585, p_wishbone_bd_ram_n22586, 
        p_wishbone_bd_ram_n22587, p_wishbone_bd_ram_n22588, 
        p_wishbone_bd_ram_n22589, p_wishbone_bd_ram_n22590, 
        p_wishbone_bd_ram_n22591, p_wishbone_bd_ram_n22592, 
        p_wishbone_bd_ram_n22593, p_wishbone_bd_ram_n22594, 
        p_wishbone_bd_ram_n22595, p_wishbone_bd_ram_n22596, 
        p_wishbone_bd_ram_n22597, p_wishbone_bd_ram_n22598, 
        p_wishbone_bd_ram_n22599, p_wishbone_bd_ram_n22600, 
        p_wishbone_bd_ram_n22601, p_wishbone_bd_ram_n22602, 
        p_wishbone_bd_ram_n22603, p_wishbone_bd_ram_n22604, 
        p_wishbone_bd_ram_n22605, p_wishbone_bd_ram_n22606, 
        p_wishbone_bd_ram_n22607, p_wishbone_bd_ram_n22608, 
        p_wishbone_bd_ram_n22609, p_wishbone_bd_ram_n22610, 
        p_wishbone_bd_ram_n22611, p_wishbone_bd_ram_n22612, 
        p_wishbone_bd_ram_n22613, p_wishbone_bd_ram_n22614, 
        p_wishbone_bd_ram_n22615, p_wishbone_bd_ram_n22616, 
        p_wishbone_bd_ram_n22617, p_wishbone_bd_ram_n22618, 
        p_wishbone_bd_ram_n22619, p_wishbone_bd_ram_n22620, 
        p_wishbone_bd_ram_n22621, p_wishbone_bd_ram_n22622, 
        p_wishbone_bd_ram_n22623, p_wishbone_bd_ram_n22624, 
        p_wishbone_bd_ram_n22625, p_wishbone_bd_ram_n22626, 
        p_wishbone_bd_ram_n22627, p_wishbone_bd_ram_n22628, 
        p_wishbone_bd_ram_n22629, p_wishbone_bd_ram_n22630, 
        p_wishbone_bd_ram_n22631, p_wishbone_bd_ram_n22632, 
        p_wishbone_bd_ram_n22633, p_wishbone_bd_ram_n22634, 
        p_wishbone_bd_ram_n22635, p_wishbone_bd_ram_n22636, 
        p_wishbone_bd_ram_n22637, p_wishbone_bd_ram_n22638, 
        p_wishbone_bd_ram_n22639, p_wishbone_bd_ram_n22640, 
        p_wishbone_bd_ram_n22641, p_wishbone_bd_ram_n22642, 
        p_wishbone_bd_ram_n22643, p_wishbone_bd_ram_n22644, 
        p_wishbone_bd_ram_n22645, p_wishbone_bd_ram_n22646, 
        p_wishbone_bd_ram_n22647, p_wishbone_bd_ram_n22648, 
        p_wishbone_bd_ram_n22649, p_wishbone_bd_ram_n22650, 
        p_wishbone_bd_ram_n22651, p_wishbone_bd_ram_n22652, 
        p_wishbone_bd_ram_n22653, p_wishbone_bd_ram_n22654, 
        p_wishbone_bd_ram_n22655, p_wishbone_bd_ram_n22656, 
        p_wishbone_bd_ram_n22657, p_wishbone_bd_ram_n22658, 
        p_wishbone_bd_ram_n22659, p_wishbone_bd_ram_n22660, 
        p_wishbone_bd_ram_n22661, p_wishbone_bd_ram_n22662, 
        p_wishbone_bd_ram_n22663, p_wishbone_bd_ram_n22664, 
        p_wishbone_bd_ram_n22665, p_wishbone_bd_ram_n22666, 
        p_wishbone_bd_ram_n22667, p_wishbone_bd_ram_n22668, 
        p_wishbone_bd_ram_n22669, p_wishbone_bd_ram_n22670, 
        p_wishbone_bd_ram_n22671, p_wishbone_bd_ram_n22672, 
        p_wishbone_bd_ram_n22673, p_wishbone_bd_ram_n22674, 
        p_wishbone_bd_ram_n22675, p_wishbone_bd_ram_n22676, 
        p_wishbone_bd_ram_n22677, p_wishbone_bd_ram_n22678, 
        p_wishbone_bd_ram_n22679, p_wishbone_bd_ram_n22680, 
        p_wishbone_bd_ram_n22681, p_wishbone_bd_ram_n22682, 
        p_wishbone_bd_ram_n22683, p_wishbone_bd_ram_n22684, 
        p_wishbone_bd_ram_n22685, p_wishbone_bd_ram_n22686, 
        p_wishbone_bd_ram_n22687, p_wishbone_bd_ram_n22688, 
        p_wishbone_bd_ram_n22689, p_wishbone_bd_ram_n22690, 
        p_wishbone_bd_ram_n22691, p_wishbone_bd_ram_n22692, 
        p_wishbone_bd_ram_n22693, p_wishbone_bd_ram_n22694, 
        p_wishbone_bd_ram_n22695, p_wishbone_bd_ram_n22696, 
        p_wishbone_bd_ram_n22697, p_wishbone_bd_ram_n22698, 
        p_wishbone_bd_ram_n22699, p_wishbone_bd_ram_n22700, 
        p_wishbone_bd_ram_n22701, p_wishbone_bd_ram_n22702, 
        p_wishbone_bd_ram_n22703, p_wishbone_bd_ram_n22704, 
        p_wishbone_bd_ram_n22705, p_wishbone_bd_ram_n22706, 
        p_wishbone_bd_ram_n22707, p_wishbone_bd_ram_n22708, 
        p_wishbone_bd_ram_n22709, p_wishbone_bd_ram_n22710, 
        p_wishbone_bd_ram_n22711, p_wishbone_bd_ram_n22712, 
        p_wishbone_bd_ram_n22713, p_wishbone_bd_ram_n22714, 
        p_wishbone_bd_ram_n22715, p_wishbone_bd_ram_n22716, 
        p_wishbone_bd_ram_n22717, p_wishbone_bd_ram_n22718, 
        p_wishbone_bd_ram_n22719, p_wishbone_bd_ram_n22720, 
        p_wishbone_bd_ram_n22721, p_wishbone_bd_ram_n22722, 
        p_wishbone_bd_ram_n22723, p_wishbone_bd_ram_n22724, 
        p_wishbone_bd_ram_n22725, p_wishbone_bd_ram_n22726, 
        p_wishbone_bd_ram_n22727, p_wishbone_bd_ram_n22728, 
        p_wishbone_bd_ram_n22729, p_wishbone_bd_ram_n22730, 
        p_wishbone_bd_ram_n22731, p_wishbone_bd_ram_n22732, 
        p_wishbone_bd_ram_n22733, p_wishbone_bd_ram_n22734, 
        p_wishbone_bd_ram_n22735, p_wishbone_bd_ram_n22736, 
        p_wishbone_bd_ram_n22737, p_wishbone_bd_ram_n22738, 
        p_wishbone_bd_ram_n22739, p_wishbone_bd_ram_n22740, 
        p_wishbone_bd_ram_n22741, p_wishbone_bd_ram_n22742, 
        p_wishbone_bd_ram_n22743, p_wishbone_bd_ram_n22744, 
        p_wishbone_bd_ram_n22745, p_wishbone_bd_ram_n22746, 
        p_wishbone_bd_ram_n22747, p_wishbone_bd_ram_n22748, 
        p_wishbone_bd_ram_n22749, p_wishbone_bd_ram_n22750, 
        p_wishbone_bd_ram_n22751, p_wishbone_bd_ram_n22752, 
        p_wishbone_bd_ram_n22753, p_wishbone_bd_ram_n22754, 
        p_wishbone_bd_ram_n22755, p_wishbone_bd_ram_n22756, 
        p_wishbone_bd_ram_n22757, p_wishbone_bd_ram_n22758, 
        p_wishbone_bd_ram_n22759, p_wishbone_bd_ram_n22760, 
        p_wishbone_bd_ram_n22761, p_wishbone_bd_ram_n22762, 
        p_wishbone_bd_ram_n22763, p_wishbone_bd_ram_n22764, 
        p_wishbone_bd_ram_n22765, p_wishbone_bd_ram_n22766, 
        p_wishbone_bd_ram_n22767, p_wishbone_bd_ram_n22768, 
        p_wishbone_bd_ram_n22769, p_wishbone_bd_ram_n22770, 
        p_wishbone_bd_ram_n22771, p_wishbone_bd_ram_n22772, 
        p_wishbone_bd_ram_n22773, p_wishbone_bd_ram_n22774, 
        p_wishbone_bd_ram_n22775, p_wishbone_bd_ram_n22776, 
        p_wishbone_bd_ram_n22777, p_wishbone_bd_ram_n22778, 
        p_wishbone_bd_ram_n22779, p_wishbone_bd_ram_n22780, 
        p_wishbone_bd_ram_n22781, p_wishbone_bd_ram_n22782, 
        p_wishbone_bd_ram_n22783, p_wishbone_bd_ram_n22784, 
        p_wishbone_bd_ram_n22785, p_wishbone_bd_ram_n22786, 
        p_wishbone_bd_ram_n22787, p_wishbone_bd_ram_n22788, 
        p_wishbone_bd_ram_n22789, p_wishbone_bd_ram_n22790, 
        p_wishbone_bd_ram_n22791, p_wishbone_bd_ram_n22792, 
        p_wishbone_bd_ram_n22793, p_wishbone_bd_ram_n22794, 
        p_wishbone_bd_ram_n22795, p_wishbone_bd_ram_n22796, 
        p_wishbone_bd_ram_n22797, p_wishbone_bd_ram_n22798, 
        p_wishbone_bd_ram_n22799, p_wishbone_bd_ram_n22800, 
        p_wishbone_bd_ram_n22801, p_wishbone_bd_ram_n22802, 
        p_wishbone_bd_ram_n22803, p_wishbone_bd_ram_n22804, 
        p_wishbone_bd_ram_n22805, p_wishbone_bd_ram_n22806, 
        p_wishbone_bd_ram_n22807, p_wishbone_bd_ram_n22808, 
        p_wishbone_bd_ram_n22809, p_wishbone_bd_ram_n22810, 
        p_wishbone_bd_ram_n22811, p_wishbone_bd_ram_n22812, 
        p_wishbone_bd_ram_n22813, p_wishbone_bd_ram_n22814, 
        p_wishbone_bd_ram_n22815, p_wishbone_bd_ram_n22816, 
        p_wishbone_bd_ram_n22817, p_wishbone_bd_ram_n22818, 
        p_wishbone_bd_ram_n22819, p_wishbone_bd_ram_n22820, 
        p_wishbone_bd_ram_n22821, p_wishbone_bd_ram_n22822, 
        p_wishbone_bd_ram_n22823, p_wishbone_bd_ram_n22824, 
        p_wishbone_bd_ram_n22825, p_wishbone_bd_ram_n22826, 
        p_wishbone_bd_ram_n22827, p_wishbone_bd_ram_n22828, 
        p_wishbone_bd_ram_n22829, p_wishbone_bd_ram_n22830, 
        p_wishbone_bd_ram_n22831, p_wishbone_bd_ram_n22832, 
        p_wishbone_bd_ram_n22833, p_wishbone_bd_ram_n22834, 
        p_wishbone_bd_ram_n22835, p_wishbone_bd_ram_n22836, 
        p_wishbone_bd_ram_n22837, p_wishbone_bd_ram_n22838, 
        p_wishbone_bd_ram_n22839, p_wishbone_bd_ram_n22840, 
        p_wishbone_bd_ram_n22841, p_wishbone_bd_ram_n22842, 
        p_wishbone_bd_ram_n22843, p_wishbone_bd_ram_n22844, 
        p_wishbone_bd_ram_n22845, p_wishbone_bd_ram_n22846, 
        p_wishbone_bd_ram_n22847, p_wishbone_bd_ram_n22848, 
        p_wishbone_bd_ram_n22849, p_wishbone_bd_ram_n22850, 
        p_wishbone_bd_ram_n22851, p_wishbone_bd_ram_n22852, 
        p_wishbone_bd_ram_n22853, p_wishbone_bd_ram_n22854, 
        p_wishbone_bd_ram_n22855, p_wishbone_bd_ram_n22856, 
        p_wishbone_bd_ram_n22857, p_wishbone_bd_ram_n22858, 
        p_wishbone_bd_ram_n22859, p_wishbone_bd_ram_n22860, 
        p_wishbone_bd_ram_n22861, p_wishbone_bd_ram_n22862, 
        p_wishbone_bd_ram_n22863, p_wishbone_bd_ram_n22864, 
        p_wishbone_bd_ram_n22865, p_wishbone_bd_ram_n22866, 
        p_wishbone_bd_ram_n22867, p_wishbone_bd_ram_n22868, 
        p_wishbone_bd_ram_n22869, p_wishbone_bd_ram_n22870, 
        p_wishbone_bd_ram_n22871, p_wishbone_bd_ram_n22872, 
        p_wishbone_bd_ram_n22873, p_wishbone_bd_ram_n22874, 
        p_wishbone_bd_ram_n22875, p_wishbone_bd_ram_n22876, 
        p_wishbone_bd_ram_n22877, p_wishbone_bd_ram_n22878, 
        p_wishbone_bd_ram_n22879, p_wishbone_bd_ram_n22880, 
        p_wishbone_bd_ram_n22881, p_wishbone_bd_ram_n22882, 
        p_wishbone_bd_ram_n22883, p_wishbone_bd_ram_n22884, 
        p_wishbone_bd_ram_n22885, p_wishbone_bd_ram_n22886, 
        p_wishbone_bd_ram_n22887, p_wishbone_bd_ram_n22888, 
        p_wishbone_bd_ram_n22889, p_wishbone_bd_ram_n22890, 
        p_wishbone_bd_ram_n22891, p_wishbone_bd_ram_n22892, 
        p_wishbone_bd_ram_n22893, p_wishbone_bd_ram_n22894, 
        p_wishbone_bd_ram_n22895, p_wishbone_bd_ram_n22896, 
        p_wishbone_bd_ram_n22897, p_wishbone_bd_ram_n22898, 
        p_wishbone_bd_ram_n22899, p_wishbone_bd_ram_n22900, 
        p_wishbone_bd_ram_n22901, p_wishbone_bd_ram_n22902, 
        p_wishbone_bd_ram_n22903, p_wishbone_bd_ram_n22904, 
        p_wishbone_bd_ram_n22905, p_wishbone_bd_ram_n22906, 
        p_wishbone_bd_ram_n22907, p_wishbone_bd_ram_n22908, 
        p_wishbone_bd_ram_n22909, p_wishbone_bd_ram_n22910, 
        p_wishbone_bd_ram_n22911, p_wishbone_bd_ram_n22912, 
        p_wishbone_bd_ram_n22913, p_wishbone_bd_ram_n22914, 
        p_wishbone_bd_ram_n22915, p_wishbone_bd_ram_n22916, 
        p_wishbone_bd_ram_n22917, p_wishbone_bd_ram_n22918, 
        p_wishbone_bd_ram_n22919, p_wishbone_bd_ram_n22920, 
        p_wishbone_bd_ram_n22921, p_wishbone_bd_ram_n22922, 
        p_wishbone_bd_ram_n22923, p_wishbone_bd_ram_n22924, 
        p_wishbone_bd_ram_n22925, p_wishbone_bd_ram_n22926, 
        p_wishbone_bd_ram_n22927, p_wishbone_bd_ram_n22928, 
        p_wishbone_bd_ram_n22929, p_wishbone_bd_ram_n22930, 
        p_wishbone_bd_ram_n22931, p_wishbone_bd_ram_n22932, 
        p_wishbone_bd_ram_n22933, p_wishbone_bd_ram_n22934, 
        p_wishbone_bd_ram_n22935, p_wishbone_bd_ram_n22936, 
        p_wishbone_bd_ram_n22937, p_wishbone_bd_ram_n22938, 
        p_wishbone_bd_ram_n22939, p_wishbone_bd_ram_n22940, 
        p_wishbone_bd_ram_n22941, p_wishbone_bd_ram_n22942, 
        p_wishbone_bd_ram_n22943, p_wishbone_bd_ram_n22944, 
        p_wishbone_bd_ram_n22945, p_wishbone_bd_ram_n22946, 
        p_wishbone_bd_ram_n22947, p_wishbone_bd_ram_n22948, 
        p_wishbone_bd_ram_n22949, p_wishbone_bd_ram_n22950, 
        p_wishbone_bd_ram_n22951, p_wishbone_bd_ram_n22952, 
        p_wishbone_bd_ram_n22953, p_wishbone_bd_ram_n22954, 
        p_wishbone_bd_ram_n22955, p_wishbone_bd_ram_n22956, 
        p_wishbone_bd_ram_n22957, p_wishbone_bd_ram_n22958, 
        p_wishbone_bd_ram_n22959, p_wishbone_bd_ram_n22960, 
        p_wishbone_bd_ram_n22961, p_wishbone_bd_ram_n22962, 
        p_wishbone_bd_ram_n22963, p_wishbone_bd_ram_n22964, 
        p_wishbone_bd_ram_n22965, p_wishbone_bd_ram_n22966, 
        p_wishbone_bd_ram_n22967, p_wishbone_bd_ram_n22968, 
        p_wishbone_bd_ram_n22969, p_wishbone_bd_ram_n22970, 
        p_wishbone_bd_ram_n22971, p_wishbone_bd_ram_n22972, 
        p_wishbone_bd_ram_n22973, p_wishbone_bd_ram_n22974, 
        p_wishbone_bd_ram_n22975, p_wishbone_bd_ram_n22976, 
        p_wishbone_bd_ram_n22977, p_wishbone_bd_ram_n22978, 
        p_wishbone_bd_ram_n22979, p_wishbone_bd_ram_n22980, 
        p_wishbone_bd_ram_n22981, p_wishbone_bd_ram_n22982, 
        p_wishbone_bd_ram_n22983, p_wishbone_bd_ram_n22984, 
        p_wishbone_bd_ram_n22985, p_wishbone_bd_ram_n22986, 
        p_wishbone_bd_ram_n22987, p_wishbone_bd_ram_n22988, 
        p_wishbone_bd_ram_n22989, p_wishbone_bd_ram_n22990, 
        p_wishbone_bd_ram_n22991, p_wishbone_bd_ram_n22992, 
        p_wishbone_bd_ram_n22993, p_wishbone_bd_ram_n22994, 
        p_wishbone_bd_ram_n22995, p_wishbone_bd_ram_n22996, 
        p_wishbone_bd_ram_n22997, p_wishbone_bd_ram_n22998, 
        p_wishbone_bd_ram_n22999, p_wishbone_bd_ram_n23000, 
        p_wishbone_bd_ram_n23001, p_wishbone_bd_ram_n23002, 
        p_wishbone_bd_ram_n23003, p_wishbone_bd_ram_n23004, 
        p_wishbone_bd_ram_n23005, p_wishbone_bd_ram_n23006, 
        p_wishbone_bd_ram_n23007, p_wishbone_bd_ram_n23008, 
        p_wishbone_bd_ram_n23009, p_wishbone_bd_ram_n23010, 
        p_wishbone_bd_ram_n23011, p_wishbone_bd_ram_n23012, 
        p_wishbone_bd_ram_n23013, p_wishbone_bd_ram_n23014, 
        p_wishbone_bd_ram_n23015, p_wishbone_bd_ram_n23016, 
        p_wishbone_bd_ram_n23017, p_wishbone_bd_ram_n23018, 
        p_wishbone_bd_ram_n23019, p_wishbone_bd_ram_n23020, 
        p_wishbone_bd_ram_n23021, p_wishbone_bd_ram_n23022, 
        p_wishbone_bd_ram_n23023, p_wishbone_bd_ram_n23024, 
        p_wishbone_bd_ram_n23025, p_wishbone_bd_ram_n23026, 
        p_wishbone_bd_ram_n23027, p_wishbone_bd_ram_n23028, 
        p_wishbone_bd_ram_n23029, p_wishbone_bd_ram_n23030, 
        p_wishbone_bd_ram_n23031, p_wishbone_bd_ram_n23032, 
        p_wishbone_bd_ram_n23033, p_wishbone_bd_ram_n23034, 
        p_wishbone_bd_ram_n23035, p_wishbone_bd_ram_n23036, 
        p_wishbone_bd_ram_n23037, p_wishbone_bd_ram_n23038, 
        p_wishbone_bd_ram_n23039, p_wishbone_bd_ram_n23040, 
        p_wishbone_bd_ram_n23041, p_wishbone_bd_ram_n23042, 
        p_wishbone_bd_ram_n23043, p_wishbone_bd_ram_n23044, 
        p_wishbone_bd_ram_n23045, p_wishbone_bd_ram_n23046, 
        p_wishbone_bd_ram_n23047, p_wishbone_bd_ram_n23048, 
        p_wishbone_bd_ram_n23049, p_wishbone_bd_ram_n23050, 
        p_wishbone_bd_ram_n23051, p_wishbone_bd_ram_n23052, 
        p_wishbone_bd_ram_n23053, p_wishbone_bd_ram_n23054, 
        p_wishbone_bd_ram_n23055, p_wishbone_bd_ram_n23056, 
        p_wishbone_bd_ram_n23057, p_wishbone_bd_ram_n23058, 
        p_wishbone_bd_ram_n23059, p_wishbone_bd_ram_n23060, 
        p_wishbone_bd_ram_n23061, p_wishbone_bd_ram_n23062, 
        p_wishbone_bd_ram_n23063, p_wishbone_bd_ram_n23064, 
        p_wishbone_bd_ram_n23065, p_wishbone_bd_ram_n23066, 
        p_wishbone_bd_ram_n23067, p_wishbone_bd_ram_n23068, 
        p_wishbone_bd_ram_n23069, p_wishbone_bd_ram_n23070, 
        p_wishbone_bd_ram_n23071, p_wishbone_bd_ram_n23072, 
        p_wishbone_bd_ram_n23073, p_wishbone_bd_ram_n23074, 
        p_wishbone_bd_ram_n23075, p_wishbone_bd_ram_n23076, 
        p_wishbone_bd_ram_n23077, p_wishbone_bd_ram_n23078, 
        p_wishbone_bd_ram_n23079, p_wishbone_bd_ram_n23080, 
        p_wishbone_bd_ram_n23081, p_wishbone_bd_ram_n23082, 
        p_wishbone_bd_ram_n23083, p_wishbone_bd_ram_n23084, 
        p_wishbone_bd_ram_n23085, p_wishbone_bd_ram_n23086, 
        p_wishbone_bd_ram_n23087, p_wishbone_bd_ram_n23088, 
        p_wishbone_bd_ram_n23089, p_wishbone_bd_ram_n23090, 
        p_wishbone_bd_ram_n23091, p_wishbone_bd_ram_n23092, 
        p_wishbone_bd_ram_n23093, p_wishbone_bd_ram_n23094, 
        p_wishbone_bd_ram_n23095, p_wishbone_bd_ram_n23096, 
        p_wishbone_bd_ram_n23097, p_wishbone_bd_ram_n23098, 
        p_wishbone_bd_ram_n23099, p_wishbone_bd_ram_n23100, 
        p_wishbone_bd_ram_n23101, p_wishbone_bd_ram_n23102, 
        p_wishbone_bd_ram_n23103, p_wishbone_bd_ram_n23104, 
        p_wishbone_bd_ram_n23105, p_wishbone_bd_ram_n23106, 
        p_wishbone_bd_ram_n23107, p_wishbone_bd_ram_n23108, 
        p_wishbone_bd_ram_n23109, p_wishbone_bd_ram_n23110, 
        p_wishbone_bd_ram_n23111, p_wishbone_bd_ram_n23112, 
        p_wishbone_bd_ram_n23113, p_wishbone_bd_ram_n23114, 
        p_wishbone_bd_ram_n23115, p_wishbone_bd_ram_n23116, 
        p_wishbone_bd_ram_n23117, p_wishbone_bd_ram_n23118, 
        p_wishbone_bd_ram_n23119, p_wishbone_bd_ram_n23120, 
        p_wishbone_bd_ram_n23121, p_wishbone_bd_ram_n23122, 
        p_wishbone_bd_ram_n23123, p_wishbone_bd_ram_n23124, 
        p_wishbone_bd_ram_n23125, p_wishbone_bd_ram_n23126, 
        p_wishbone_bd_ram_n23127, p_wishbone_bd_ram_n23128, 
        p_wishbone_bd_ram_n23129, p_wishbone_bd_ram_n23130, 
        p_wishbone_bd_ram_n23131, p_wishbone_bd_ram_n23132, 
        p_wishbone_bd_ram_n23133, p_wishbone_bd_ram_n23134, 
        p_wishbone_bd_ram_n23135, p_wishbone_bd_ram_n23136, 
        p_wishbone_bd_ram_n23137, p_wishbone_bd_ram_n23138, 
        p_wishbone_bd_ram_n23139, p_wishbone_bd_ram_n23140, 
        p_wishbone_bd_ram_n23141, p_wishbone_bd_ram_n23142, 
        p_wishbone_bd_ram_n23143, p_wishbone_bd_ram_n23144, 
        p_wishbone_bd_ram_n23145, p_wishbone_bd_ram_n23146, 
        p_wishbone_bd_ram_n23147, p_wishbone_bd_ram_n23148, 
        p_wishbone_bd_ram_n23149, p_wishbone_bd_ram_n23150, 
        p_wishbone_bd_ram_n23151, p_wishbone_bd_ram_n23152, 
        p_wishbone_bd_ram_n23153, p_wishbone_bd_ram_n23154, 
        p_wishbone_bd_ram_n23155, p_wishbone_bd_ram_n23156, 
        p_wishbone_bd_ram_n23157, p_wishbone_bd_ram_n23158, 
        p_wishbone_bd_ram_n23159, p_wishbone_bd_ram_n23160, 
        p_wishbone_bd_ram_n23161, p_wishbone_bd_ram_n23162, 
        p_wishbone_bd_ram_n23163, p_wishbone_bd_ram_n23164, 
        p_wishbone_bd_ram_n23165, p_wishbone_bd_ram_n23166, 
        p_wishbone_bd_ram_n23167, p_wishbone_bd_ram_n23168, 
        p_wishbone_bd_ram_n23169, p_wishbone_bd_ram_n23170, 
        p_wishbone_bd_ram_n23171, p_wishbone_bd_ram_n23172, 
        p_wishbone_bd_ram_n23173, p_wishbone_bd_ram_n23174, 
        p_wishbone_bd_ram_n23175, p_wishbone_bd_ram_n23176, 
        p_wishbone_bd_ram_n23177, p_wishbone_bd_ram_n23178, 
        p_wishbone_bd_ram_n23179, p_wishbone_bd_ram_n23180, 
        p_wishbone_bd_ram_n23181, p_wishbone_bd_ram_n23182, 
        p_wishbone_bd_ram_n23183, p_wishbone_bd_ram_n23184, 
        p_wishbone_bd_ram_n23185, p_wishbone_bd_ram_n23186, 
        p_wishbone_bd_ram_n23187, p_wishbone_bd_ram_n23188, 
        p_wishbone_bd_ram_n23189, p_wishbone_bd_ram_n23190, 
        p_wishbone_bd_ram_n23191, p_wishbone_bd_ram_n23192, 
        p_wishbone_bd_ram_n23193, p_wishbone_bd_ram_n23194, 
        p_wishbone_bd_ram_n23195, p_wishbone_bd_ram_n23196, 
        p_wishbone_bd_ram_n23197, p_wishbone_bd_ram_n23198, 
        p_wishbone_bd_ram_n23199, p_wishbone_bd_ram_n23200, 
        p_wishbone_bd_ram_n23201, p_wishbone_bd_ram_n23202, 
        p_wishbone_bd_ram_n23203, p_wishbone_bd_ram_n23204, 
        p_wishbone_bd_ram_n23205, p_wishbone_bd_ram_n23206, 
        p_wishbone_bd_ram_n23207, p_wishbone_bd_ram_n23208, 
        p_wishbone_bd_ram_n23209, p_wishbone_bd_ram_n23210, 
        p_wishbone_bd_ram_n23211, p_wishbone_bd_ram_n23212, 
        p_wishbone_bd_ram_n23213, p_wishbone_bd_ram_n23214, 
        p_wishbone_bd_ram_n23215, p_wishbone_bd_ram_n23216, 
        p_wishbone_bd_ram_n23217, p_wishbone_bd_ram_n23218, 
        p_wishbone_bd_ram_n23219, p_wishbone_bd_ram_n23220, 
        p_wishbone_bd_ram_n23221, p_wishbone_bd_ram_n23222, 
        p_wishbone_bd_ram_n23223, p_wishbone_bd_ram_n23224, 
        p_wishbone_bd_ram_n23225, p_wishbone_bd_ram_n23226, 
        p_wishbone_bd_ram_n23227, p_wishbone_bd_ram_n23228, 
        p_wishbone_bd_ram_n23229, p_wishbone_bd_ram_n23230, 
        p_wishbone_bd_ram_n23231, p_wishbone_bd_ram_n23232, 
        p_wishbone_bd_ram_n23233, p_wishbone_bd_ram_n23234, 
        p_wishbone_bd_ram_n23235, p_wishbone_bd_ram_n23236, 
        p_wishbone_bd_ram_n23237, p_wishbone_bd_ram_n23238, 
        p_wishbone_bd_ram_n23239, p_wishbone_bd_ram_n23240, 
        p_wishbone_bd_ram_n23241, p_wishbone_bd_ram_n23242, 
        p_wishbone_bd_ram_n23243, p_wishbone_bd_ram_n23244, 
        p_wishbone_bd_ram_n23245, p_wishbone_bd_ram_n23246, 
        p_wishbone_bd_ram_n23247, p_wishbone_bd_ram_n23248, 
        p_wishbone_bd_ram_n23249, p_wishbone_bd_ram_n23250, 
        p_wishbone_bd_ram_n23251, p_wishbone_bd_ram_n23252, 
        p_wishbone_bd_ram_n23253, p_wishbone_bd_ram_n23254, 
        p_wishbone_bd_ram_n23255, p_wishbone_bd_ram_n23256, 
        p_wishbone_bd_ram_n23257, p_wishbone_bd_ram_n23258, 
        p_wishbone_bd_ram_n23259, p_wishbone_bd_ram_n23260, 
        p_wishbone_bd_ram_n23261, p_wishbone_bd_ram_n23262, 
        p_wishbone_bd_ram_n23263, p_wishbone_bd_ram_n23264, 
        p_wishbone_bd_ram_n23265, p_wishbone_bd_ram_n23266, 
        p_wishbone_bd_ram_n23267, p_wishbone_bd_ram_n23268, 
        p_wishbone_bd_ram_n23269, p_wishbone_bd_ram_n23270, 
        p_wishbone_bd_ram_n23271, p_wishbone_bd_ram_n23272, 
        p_wishbone_bd_ram_n23273, p_wishbone_bd_ram_n23274, 
        p_wishbone_bd_ram_n23275, p_wishbone_bd_ram_n23276, 
        p_wishbone_bd_ram_n23277, p_wishbone_bd_ram_n23278, 
        p_wishbone_bd_ram_n23279, p_wishbone_bd_ram_n23280, 
        p_wishbone_bd_ram_n23281, p_wishbone_bd_ram_n23282, 
        p_wishbone_bd_ram_n23283, p_wishbone_bd_ram_n23284, 
        p_wishbone_bd_ram_n23285, p_wishbone_bd_ram_n23286, 
        p_wishbone_bd_ram_n23287, p_wishbone_bd_ram_n23288, 
        p_wishbone_bd_ram_n23289, p_wishbone_bd_ram_n23290, 
        p_wishbone_bd_ram_n23291, p_wishbone_bd_ram_n23292, 
        p_wishbone_bd_ram_n23293, p_wishbone_bd_ram_n23294, 
        p_wishbone_bd_ram_n23295, p_wishbone_bd_ram_n23296, 
        p_wishbone_bd_ram_n23297, p_wishbone_bd_ram_n23298, 
        p_wishbone_bd_ram_n23299, p_wishbone_bd_ram_n23300, 
        p_wishbone_bd_ram_n23301, p_wishbone_bd_ram_n23302, 
        p_wishbone_bd_ram_n23303, p_wishbone_bd_ram_n23304, 
        p_wishbone_bd_ram_n23305, p_wishbone_bd_ram_n23306, 
        p_wishbone_bd_ram_n23307, p_wishbone_bd_ram_n23308, 
        p_wishbone_bd_ram_n23309, p_wishbone_bd_ram_n23310, 
        p_wishbone_bd_ram_n23311, p_wishbone_bd_ram_n23312, 
        p_wishbone_bd_ram_n23313, p_wishbone_bd_ram_n23314, 
        p_wishbone_bd_ram_n23315, p_wishbone_bd_ram_n23316, 
        p_wishbone_bd_ram_n23317, p_wishbone_bd_ram_n23318, 
        p_wishbone_bd_ram_n23319, p_wishbone_bd_ram_n23320, 
        p_wishbone_bd_ram_n23321, p_wishbone_bd_ram_n23322, 
        p_wishbone_bd_ram_n23323, p_wishbone_bd_ram_n23324, 
        p_wishbone_bd_ram_n23325, p_wishbone_bd_ram_n23326, 
        p_wishbone_bd_ram_n23327, p_wishbone_bd_ram_n23328, 
        p_wishbone_bd_ram_n23329, p_wishbone_bd_ram_n23330, 
        p_wishbone_bd_ram_n23331, p_wishbone_bd_ram_n23332, 
        p_wishbone_bd_ram_n23333, p_wishbone_bd_ram_n23334, 
        p_wishbone_bd_ram_n23335, p_wishbone_bd_ram_n23336, 
        p_wishbone_bd_ram_n23337, p_wishbone_bd_ram_n23338, 
        p_wishbone_bd_ram_n23339, p_wishbone_bd_ram_n23340, 
        p_wishbone_bd_ram_n23341, p_wishbone_bd_ram_n23342, 
        p_wishbone_bd_ram_n23343, p_wishbone_bd_ram_n23344, 
        p_wishbone_bd_ram_n23345, p_wishbone_bd_ram_n23346, 
        p_wishbone_bd_ram_n23347, p_wishbone_bd_ram_n23348, 
        p_wishbone_bd_ram_n23349, p_wishbone_bd_ram_n23350, 
        p_wishbone_bd_ram_n23351, p_wishbone_bd_ram_n23352, 
        p_wishbone_bd_ram_n23353, p_wishbone_bd_ram_n23354, 
        p_wishbone_bd_ram_n23355, p_wishbone_bd_ram_n23356, 
        p_wishbone_bd_ram_n23357, p_wishbone_bd_ram_n23358, 
        p_wishbone_bd_ram_n23359, p_wishbone_bd_ram_n23360, 
        p_wishbone_bd_ram_n23361, p_wishbone_bd_ram_n23362, 
        p_wishbone_bd_ram_n23363, p_wishbone_bd_ram_n23364, 
        p_wishbone_bd_ram_n23365, p_wishbone_bd_ram_n23366, 
        p_wishbone_bd_ram_n23367, p_wishbone_bd_ram_n23368, 
        p_wishbone_bd_ram_n23369, p_wishbone_bd_ram_n23370, 
        p_wishbone_bd_ram_n23371, p_wishbone_bd_ram_n23372, 
        p_wishbone_bd_ram_n23373, p_wishbone_bd_ram_n23374, 
        p_wishbone_bd_ram_n23375, p_wishbone_bd_ram_n23376, 
        p_wishbone_bd_ram_n23377, p_wishbone_bd_ram_n23378, 
        p_wishbone_bd_ram_n23379, p_wishbone_bd_ram_n23380, 
        p_wishbone_bd_ram_n23381, p_wishbone_bd_ram_n23382, 
        p_wishbone_bd_ram_n23383, p_wishbone_bd_ram_n23384, 
        p_wishbone_bd_ram_n23385, p_wishbone_bd_ram_n23386, 
        p_wishbone_bd_ram_n23387, p_wishbone_bd_ram_n23388, 
        p_wishbone_bd_ram_n23389, p_wishbone_bd_ram_n23390, 
        p_wishbone_bd_ram_n23391, p_wishbone_bd_ram_n23392, 
        p_wishbone_bd_ram_n23393, p_wishbone_bd_ram_n23394, 
        p_wishbone_bd_ram_n23395, p_wishbone_bd_ram_n23396, 
        p_wishbone_bd_ram_n23397, p_wishbone_bd_ram_n23398, 
        p_wishbone_bd_ram_n23399, p_wishbone_bd_ram_n23400, 
        p_wishbone_bd_ram_n23401, p_wishbone_bd_ram_n23402, 
        p_wishbone_bd_ram_n23403, p_wishbone_bd_ram_n23404, 
        p_wishbone_bd_ram_n23405, p_wishbone_bd_ram_n23406, 
        p_wishbone_bd_ram_n23407, p_wishbone_bd_ram_n23408, 
        p_wishbone_bd_ram_n23409, p_wishbone_bd_ram_n23410, 
        p_wishbone_bd_ram_n23411, p_wishbone_bd_ram_n23412, 
        p_wishbone_bd_ram_n23413, p_wishbone_bd_ram_n23414, 
        p_wishbone_bd_ram_n23415, p_wishbone_bd_ram_n23416, 
        p_wishbone_bd_ram_n23417, p_wishbone_bd_ram_n23418, 
        p_wishbone_bd_ram_n23419, p_wishbone_bd_ram_n23420, 
        p_wishbone_bd_ram_n23421, p_wishbone_bd_ram_n23422, 
        p_wishbone_bd_ram_n23423, p_wishbone_bd_ram_n23424, 
        p_wishbone_bd_ram_n23425, p_wishbone_bd_ram_n23426, 
        p_wishbone_bd_ram_n23427, p_wishbone_bd_ram_n23428, 
        p_wishbone_bd_ram_n23429, p_wishbone_bd_ram_n23430, 
        p_wishbone_bd_ram_n23431, p_wishbone_bd_ram_n23432, 
        p_wishbone_bd_ram_n23433, p_wishbone_bd_ram_n23434, 
        p_wishbone_bd_ram_n23435, p_wishbone_bd_ram_n23436, 
        p_wishbone_bd_ram_n23437, p_wishbone_bd_ram_n23438, 
        p_wishbone_bd_ram_n23439, p_wishbone_bd_ram_n23440, 
        p_wishbone_bd_ram_n23441, p_wishbone_bd_ram_n23442, 
        p_wishbone_bd_ram_n23443, p_wishbone_bd_ram_n23444, 
        p_wishbone_bd_ram_n23445, p_wishbone_bd_ram_n23446, 
        p_wishbone_bd_ram_n23447, p_wishbone_bd_ram_n23448, 
        p_wishbone_bd_ram_n23449, p_wishbone_bd_ram_n23450, 
        p_wishbone_bd_ram_n23451, p_wishbone_bd_ram_n23452, 
        p_wishbone_bd_ram_n23453, p_wishbone_bd_ram_n23454, 
        p_wishbone_bd_ram_n23455, p_wishbone_bd_ram_n23456, 
        p_wishbone_bd_ram_n23457, p_wishbone_bd_ram_n23458, 
        p_wishbone_bd_ram_n23459, p_wishbone_bd_ram_n23460, 
        p_wishbone_bd_ram_n23461, p_wishbone_bd_ram_n23462, 
        p_wishbone_bd_ram_n23463, p_wishbone_bd_ram_n23464, 
        p_wishbone_bd_ram_n23465, p_wishbone_bd_ram_n23466, 
        p_wishbone_bd_ram_n23467, p_wishbone_bd_ram_n23468, 
        p_wishbone_bd_ram_n23469, p_wishbone_bd_ram_n23470, 
        p_wishbone_bd_ram_n23471, p_wishbone_bd_ram_n23472, 
        p_wishbone_bd_ram_n23473, p_wishbone_bd_ram_n23474, 
        p_wishbone_bd_ram_n23475, p_wishbone_bd_ram_n23476, 
        p_wishbone_bd_ram_n23477, p_wishbone_bd_ram_n23478, 
        p_wishbone_bd_ram_n23479, p_wishbone_bd_ram_n23480, 
        p_wishbone_bd_ram_n23481, p_wishbone_bd_ram_n23482, 
        p_wishbone_bd_ram_n23483, p_wishbone_bd_ram_n23484, 
        p_wishbone_bd_ram_n23485, p_wishbone_bd_ram_n23486, 
        p_wishbone_bd_ram_n23487, p_wishbone_bd_ram_n23488, 
        p_wishbone_bd_ram_n23489, p_wishbone_bd_ram_n23490, 
        p_wishbone_bd_ram_n23491, p_wishbone_bd_ram_n23492, 
        p_wishbone_bd_ram_n23493, p_wishbone_bd_ram_n23494, 
        p_wishbone_bd_ram_n23495, p_wishbone_bd_ram_n23496, 
        p_wishbone_bd_ram_n23497, p_wishbone_bd_ram_n23498, 
        p_wishbone_bd_ram_n23499, p_wishbone_bd_ram_n23500, 
        p_wishbone_bd_ram_n23501, p_wishbone_bd_ram_n23502, 
        p_wishbone_bd_ram_n23503, p_wishbone_bd_ram_n23504, 
        p_wishbone_bd_ram_n23505, p_wishbone_bd_ram_n23506, 
        p_wishbone_bd_ram_n23507, p_wishbone_bd_ram_n23508, 
        p_wishbone_bd_ram_n23509, p_wishbone_bd_ram_n23510, 
        p_wishbone_bd_ram_n23511, p_wishbone_bd_ram_n23512, 
        p_wishbone_bd_ram_n23513, p_wishbone_bd_ram_n23514, 
        p_wishbone_bd_ram_n23515, p_wishbone_bd_ram_n23516, 
        p_wishbone_bd_ram_n23517, p_wishbone_bd_ram_n23518, 
        p_wishbone_bd_ram_n23519, p_wishbone_bd_ram_n23520, 
        p_wishbone_bd_ram_n23521, p_wishbone_bd_ram_n23522, 
        p_wishbone_bd_ram_n23523, p_wishbone_bd_ram_n23524, 
        p_wishbone_bd_ram_n23525, p_wishbone_bd_ram_n23526, 
        p_wishbone_bd_ram_n23527, p_wishbone_bd_ram_n23528, 
        p_wishbone_bd_ram_n23529, p_wishbone_bd_ram_n23530, 
        p_wishbone_bd_ram_n23531, p_wishbone_bd_ram_n23532, 
        p_wishbone_bd_ram_n23533, p_wishbone_bd_ram_n23534, 
        p_wishbone_bd_ram_n23535, p_wishbone_bd_ram_n23536, 
        p_wishbone_bd_ram_n23537, p_wishbone_bd_ram_n23538, 
        p_wishbone_bd_ram_n23539, p_wishbone_bd_ram_n23540, 
        p_wishbone_bd_ram_n23541, p_wishbone_bd_ram_n23542, 
        p_wishbone_bd_ram_n23543, p_wishbone_bd_ram_n23544, 
        p_wishbone_bd_ram_n23545, p_wishbone_bd_ram_n23546, 
        p_wishbone_bd_ram_n23547, p_wishbone_bd_ram_n23548, 
        p_wishbone_bd_ram_n23549, p_wishbone_bd_ram_n23550, 
        p_wishbone_bd_ram_n23551, p_wishbone_bd_ram_n23552, 
        p_wishbone_bd_ram_n23553, p_wishbone_bd_ram_n23554, 
        p_wishbone_bd_ram_n23555, p_wishbone_bd_ram_n23556, 
        p_wishbone_bd_ram_n23557, p_wishbone_bd_ram_n23558, 
        p_wishbone_bd_ram_n23559, p_wishbone_bd_ram_n23560, 
        p_wishbone_bd_ram_n23561, p_wishbone_bd_ram_n23562, 
        p_wishbone_bd_ram_n23563, p_wishbone_bd_ram_n23564, 
        p_wishbone_bd_ram_n23565, p_wishbone_bd_ram_n23566, 
        p_wishbone_bd_ram_n23567, p_wishbone_bd_ram_n23568, 
        p_wishbone_bd_ram_n23569, p_wishbone_bd_ram_n23570, 
        p_wishbone_bd_ram_n23571, p_wishbone_bd_ram_n23572, 
        p_wishbone_bd_ram_n23573, p_wishbone_bd_ram_n23574, 
        p_wishbone_bd_ram_n23575, p_wishbone_bd_ram_n23576, 
        p_wishbone_bd_ram_n23577, p_wishbone_bd_ram_n23578, 
        p_wishbone_bd_ram_n23579, p_wishbone_bd_ram_n23580, 
        p_wishbone_bd_ram_n23581, p_wishbone_bd_ram_n23582, 
        p_wishbone_bd_ram_n23583, p_wishbone_bd_ram_n23584, 
        p_wishbone_bd_ram_n23585, p_wishbone_bd_ram_n23586, 
        p_wishbone_bd_ram_n23587, p_wishbone_bd_ram_n23588, 
        p_wishbone_bd_ram_n23589, p_wishbone_bd_ram_n23590, 
        p_wishbone_bd_ram_n23591, p_wishbone_bd_ram_n23592, 
        p_wishbone_bd_ram_n23593, p_wishbone_bd_ram_n23594, 
        p_wishbone_bd_ram_n23595, p_wishbone_bd_ram_n23596, 
        p_wishbone_bd_ram_n23597, p_wishbone_bd_ram_n23598, 
        p_wishbone_bd_ram_n23599, p_wishbone_bd_ram_n23600, 
        p_wishbone_bd_ram_n23601, p_wishbone_bd_ram_n23602, 
        p_wishbone_bd_ram_n23603, p_wishbone_bd_ram_n23604, 
        p_wishbone_bd_ram_n23605, p_wishbone_bd_ram_n23606, 
        p_wishbone_bd_ram_n23607, p_wishbone_bd_ram_n23608, 
        p_wishbone_bd_ram_n23609, p_wishbone_bd_ram_n23610, 
        p_wishbone_bd_ram_n23611, p_wishbone_bd_ram_n23612, 
        p_wishbone_bd_ram_n23613, p_wishbone_bd_ram_n23614, 
        p_wishbone_bd_ram_n23615, p_wishbone_bd_ram_n23616, 
        p_wishbone_bd_ram_n23617, p_wishbone_bd_ram_n23618, 
        p_wishbone_bd_ram_n23619, p_wishbone_bd_ram_n23620, 
        p_wishbone_bd_ram_n23621, p_wishbone_bd_ram_n23622, 
        p_wishbone_bd_ram_n23623, p_wishbone_bd_ram_n23624, 
        p_wishbone_bd_ram_n23625, p_wishbone_bd_ram_n23626, 
        p_wishbone_bd_ram_n23627, p_wishbone_bd_ram_n23628, 
        p_wishbone_bd_ram_n23629, p_wishbone_bd_ram_n23630, 
        p_wishbone_bd_ram_n23631, p_wishbone_bd_ram_n23632, 
        p_wishbone_bd_ram_n23633, p_wishbone_bd_ram_n23634, 
        p_wishbone_bd_ram_n23635, p_wishbone_bd_ram_n23636, 
        p_wishbone_bd_ram_n23637, p_wishbone_bd_ram_n23638, 
        p_wishbone_bd_ram_n23639, p_wishbone_bd_ram_n23640, 
        p_wishbone_bd_ram_n23641, p_wishbone_bd_ram_n23642, 
        p_wishbone_bd_ram_n23643, p_wishbone_bd_ram_n23644, 
        p_wishbone_bd_ram_n23645, p_wishbone_bd_ram_n23646, 
        p_wishbone_bd_ram_n23647, p_wishbone_bd_ram_n23648, 
        p_wishbone_bd_ram_n23649, p_wishbone_bd_ram_n23650, 
        p_wishbone_bd_ram_n23651, p_wishbone_bd_ram_n23652, 
        p_wishbone_bd_ram_n23653, p_wishbone_bd_ram_n23654, 
        p_wishbone_bd_ram_n23655, p_wishbone_bd_ram_n23656, 
        p_wishbone_bd_ram_n23657, p_wishbone_bd_ram_n23658, 
        p_wishbone_bd_ram_n23659, p_wishbone_bd_ram_n23660, 
        p_wishbone_bd_ram_n23661, p_wishbone_bd_ram_n23662, 
        p_wishbone_bd_ram_n23663, p_wishbone_bd_ram_n23664, 
        p_wishbone_bd_ram_n23665, p_wishbone_bd_ram_n23666, 
        p_wishbone_bd_ram_n23667, p_wishbone_bd_ram_n23668, 
        p_wishbone_bd_ram_n23669, p_wishbone_bd_ram_n23670, 
        p_wishbone_bd_ram_n23671, p_wishbone_bd_ram_n23672, 
        p_wishbone_bd_ram_n23673, p_wishbone_bd_ram_n23674, 
        p_wishbone_bd_ram_n23675, p_wishbone_bd_ram_n23676, 
        p_wishbone_bd_ram_n23677, p_wishbone_bd_ram_n23678, 
        p_wishbone_bd_ram_n23679, p_wishbone_bd_ram_n23680, 
        p_wishbone_bd_ram_n23681, p_wishbone_bd_ram_n23682, 
        p_wishbone_bd_ram_n23683, p_wishbone_bd_ram_n23684, 
        p_wishbone_bd_ram_n23685, p_wishbone_bd_ram_n23686, 
        p_wishbone_bd_ram_n23687, p_wishbone_bd_ram_n23688, 
        p_wishbone_bd_ram_n23689, p_wishbone_bd_ram_n23690, 
        p_wishbone_bd_ram_n23691, p_wishbone_bd_ram_n23692, 
        p_wishbone_bd_ram_n23693, p_wishbone_bd_ram_n23694, 
        p_wishbone_bd_ram_n23695, p_wishbone_bd_ram_n23696, 
        p_wishbone_bd_ram_n23697, p_wishbone_bd_ram_n23698, 
        p_wishbone_bd_ram_n23699, p_wishbone_bd_ram_n23700, 
        p_wishbone_bd_ram_n23701, p_wishbone_bd_ram_n23702, 
        p_wishbone_bd_ram_n23703, p_wishbone_bd_ram_n23704, 
        p_wishbone_bd_ram_n23705, p_wishbone_bd_ram_n23706, 
        p_wishbone_bd_ram_n23707, p_wishbone_bd_ram_n23708, 
        p_wishbone_bd_ram_n23709, p_wishbone_bd_ram_n23710, 
        p_wishbone_bd_ram_n23711, p_wishbone_bd_ram_n23712, 
        p_wishbone_bd_ram_n23713, p_wishbone_bd_ram_n23714, 
        p_wishbone_bd_ram_n23715, p_wishbone_bd_ram_n23716, 
        p_wishbone_bd_ram_n23717, p_wishbone_bd_ram_n23718, 
        p_wishbone_bd_ram_n23719, p_wishbone_bd_ram_n23720, 
        p_wishbone_bd_ram_n23721, p_wishbone_bd_ram_n23722, 
        p_wishbone_bd_ram_n23723, p_wishbone_bd_ram_n23724, 
        p_wishbone_bd_ram_n23725, p_wishbone_bd_ram_n23726, 
        p_wishbone_bd_ram_n23727, p_wishbone_bd_ram_n23728, 
        p_wishbone_bd_ram_n23729, p_wishbone_bd_ram_n23730, 
        p_wishbone_bd_ram_n23731, p_wishbone_bd_ram_n23732, 
        p_wishbone_bd_ram_n23733, p_wishbone_bd_ram_n23734, 
        p_wishbone_bd_ram_n23735, p_wishbone_bd_ram_n23736, 
        p_wishbone_bd_ram_n23737, p_wishbone_bd_ram_n23738, 
        p_wishbone_bd_ram_n23739, p_wishbone_bd_ram_n23740, 
        p_wishbone_bd_ram_n23741, p_wishbone_bd_ram_n23742, 
        p_wishbone_bd_ram_n23743, p_wishbone_bd_ram_n23744, 
        p_wishbone_bd_ram_n23745, p_wishbone_bd_ram_n23746, 
        p_wishbone_bd_ram_n23747, p_wishbone_bd_ram_n23748, 
        p_wishbone_bd_ram_n23749, p_wishbone_bd_ram_n23750, 
        p_wishbone_bd_ram_n23751, p_wishbone_bd_ram_n23752, 
        p_wishbone_bd_ram_n23753, p_wishbone_bd_ram_n23754, 
        p_wishbone_bd_ram_n23755, p_wishbone_bd_ram_n23756, 
        p_wishbone_bd_ram_n23757, p_wishbone_bd_ram_n23758, 
        p_wishbone_bd_ram_n23759, p_wishbone_bd_ram_n23760, 
        p_wishbone_bd_ram_n23761, p_wishbone_bd_ram_n23762, 
        p_wishbone_bd_ram_n23763, p_wishbone_bd_ram_n23764, 
        p_wishbone_bd_ram_n23765, p_wishbone_bd_ram_n23766, 
        p_wishbone_bd_ram_n23767, p_wishbone_bd_ram_n23768, 
        p_wishbone_bd_ram_n23769, p_wishbone_bd_ram_n23770, 
        p_wishbone_bd_ram_n23771, p_wishbone_bd_ram_n23772, 
        p_wishbone_bd_ram_n23773, p_wishbone_bd_ram_n23774, 
        p_wishbone_bd_ram_n23775, p_wishbone_bd_ram_n23776, 
        p_wishbone_bd_ram_n23777, p_wishbone_bd_ram_n23778, 
        p_wishbone_bd_ram_n23779, p_wishbone_bd_ram_n23780, 
        p_wishbone_bd_ram_n23781, p_wishbone_bd_ram_n23782, 
        p_wishbone_bd_ram_n23783, p_wishbone_bd_ram_n23784, 
        p_wishbone_bd_ram_n23785, p_wishbone_bd_ram_n23786, 
        p_wishbone_bd_ram_n23787, p_wishbone_bd_ram_n23788, 
        p_wishbone_bd_ram_n23789, p_wishbone_bd_ram_n23790, 
        p_wishbone_bd_ram_n23791, p_wishbone_bd_ram_n23792, 
        p_wishbone_bd_ram_n23793, p_wishbone_bd_ram_n23794, 
        p_wishbone_bd_ram_n23795, p_wishbone_bd_ram_n23796, 
        p_wishbone_bd_ram_n23797, p_wishbone_bd_ram_n23798, 
        p_wishbone_bd_ram_n23799, p_wishbone_bd_ram_n23800, 
        p_wishbone_bd_ram_n23801, p_wishbone_bd_ram_n23802, 
        p_wishbone_bd_ram_n23803, p_wishbone_bd_ram_n23804, 
        p_wishbone_bd_ram_n23805, p_wishbone_bd_ram_n23806, 
        p_wishbone_bd_ram_n23807, p_wishbone_bd_ram_n23808, 
        p_wishbone_bd_ram_n23809, p_wishbone_bd_ram_n23810, 
        p_wishbone_bd_ram_n23811, p_wishbone_bd_ram_n23812, 
        p_wishbone_bd_ram_n23813, p_wishbone_bd_ram_n23814, 
        p_wishbone_bd_ram_n23815, p_wishbone_bd_ram_n23816, 
        p_wishbone_bd_ram_n23817, p_wishbone_bd_ram_n23818, 
        p_wishbone_bd_ram_n23819, p_wishbone_bd_ram_n23820, 
        p_wishbone_bd_ram_n23821, p_wishbone_bd_ram_n23822, 
        p_wishbone_bd_ram_n23823, p_wishbone_bd_ram_n23824, 
        p_wishbone_bd_ram_n23825, p_wishbone_bd_ram_n23826, 
        p_wishbone_bd_ram_n23827, p_wishbone_bd_ram_n23828, 
        p_wishbone_bd_ram_n23829, p_wishbone_bd_ram_n23830, 
        p_wishbone_bd_ram_n23831, p_wishbone_bd_ram_n23832, 
        p_wishbone_bd_ram_n23833, p_wishbone_bd_ram_n23834, 
        p_wishbone_bd_ram_n23835, p_wishbone_bd_ram_n23836, 
        p_wishbone_bd_ram_n23837, p_wishbone_bd_ram_n23838, 
        p_wishbone_bd_ram_n23839, p_wishbone_bd_ram_n23840, 
        p_wishbone_bd_ram_n23841, p_wishbone_bd_ram_n23842, 
        p_wishbone_bd_ram_n23843, p_wishbone_bd_ram_n23844, 
        p_wishbone_bd_ram_n23845, p_wishbone_bd_ram_n23846, 
        p_wishbone_bd_ram_n23847, p_wishbone_bd_ram_n23848, 
        p_wishbone_bd_ram_n23849, p_wishbone_bd_ram_n23850, 
        p_wishbone_bd_ram_n23851, p_wishbone_bd_ram_n23852, 
        p_wishbone_bd_ram_n23853, p_wishbone_bd_ram_n23854, 
        p_wishbone_bd_ram_n23855, p_wishbone_bd_ram_n23856, 
        p_wishbone_bd_ram_n23857, p_wishbone_bd_ram_n23858, 
        p_wishbone_bd_ram_n23859, p_wishbone_bd_ram_n23860, 
        p_wishbone_bd_ram_n23861, p_wishbone_bd_ram_n23862, 
        p_wishbone_bd_ram_n23863, p_wishbone_bd_ram_n23864, 
        p_wishbone_bd_ram_n23865, p_wishbone_bd_ram_n23866, 
        p_wishbone_bd_ram_n23867, p_wishbone_bd_ram_n23868, 
        p_wishbone_bd_ram_n23869, p_wishbone_bd_ram_n23870, 
        p_wishbone_bd_ram_n23871, p_wishbone_bd_ram_n23872, 
        p_wishbone_bd_ram_n23873, p_wishbone_bd_ram_n23874, 
        p_wishbone_bd_ram_n23875, p_wishbone_bd_ram_n23876, 
        p_wishbone_bd_ram_n23877, p_wishbone_bd_ram_n23878, 
        p_wishbone_bd_ram_n23879, p_wishbone_bd_ram_n23880, 
        p_wishbone_bd_ram_n23881, p_wishbone_bd_ram_n23882, 
        p_wishbone_bd_ram_n23883, p_wishbone_bd_ram_n23884, 
        p_wishbone_bd_ram_n23885, p_wishbone_bd_ram_n23886, 
        p_wishbone_bd_ram_n23887, p_wishbone_bd_ram_n23888, 
        p_wishbone_bd_ram_n23889, p_wishbone_bd_ram_n23890, 
        p_wishbone_bd_ram_n23891, p_wishbone_bd_ram_n23892, 
        p_wishbone_bd_ram_n23893, p_wishbone_bd_ram_n23894, 
        p_wishbone_bd_ram_n23895, p_wishbone_bd_ram_n23896, 
        p_wishbone_bd_ram_n23897, p_wishbone_bd_ram_n23898, 
        p_wishbone_bd_ram_n23899, p_wishbone_bd_ram_n23900, 
        p_wishbone_bd_ram_n23901, p_wishbone_bd_ram_n23902, 
        p_wishbone_bd_ram_n23903, p_wishbone_bd_ram_n23904, 
        p_wishbone_bd_ram_n23905, p_wishbone_bd_ram_n23906, 
        p_wishbone_bd_ram_n23907, p_wishbone_bd_ram_n23908, 
        p_wishbone_bd_ram_n23909, p_wishbone_bd_ram_n23910, 
        p_wishbone_bd_ram_n23911, p_wishbone_bd_ram_n23912, 
        p_wishbone_bd_ram_n23913, p_wishbone_bd_ram_n23914, 
        p_wishbone_bd_ram_n23915, p_wishbone_bd_ram_n23916, 
        p_wishbone_bd_ram_n23917, p_wishbone_bd_ram_n23918, 
        p_wishbone_bd_ram_n23919, p_wishbone_bd_ram_n23920, 
        p_wishbone_bd_ram_n23921, p_wishbone_bd_ram_n23922, 
        p_wishbone_bd_ram_n23923, p_wishbone_bd_ram_n23924, 
        p_wishbone_bd_ram_n23925, p_wishbone_bd_ram_n23926, 
        p_wishbone_bd_ram_n23927, p_wishbone_bd_ram_n23928, 
        p_wishbone_bd_ram_n23929, p_wishbone_bd_ram_n23930, 
        p_wishbone_bd_ram_n23931, p_wishbone_bd_ram_n23932, 
        p_wishbone_bd_ram_n23933, p_wishbone_bd_ram_n23934, 
        p_wishbone_bd_ram_n23935, p_wishbone_bd_ram_n23936, 
        p_wishbone_bd_ram_n23937, p_wishbone_bd_ram_n23938, 
        p_wishbone_bd_ram_n23939, p_wishbone_bd_ram_n23940, 
        p_wishbone_bd_ram_n23941, p_wishbone_bd_ram_n23942, 
        p_wishbone_bd_ram_n23943, p_wishbone_bd_ram_n23944, 
        p_wishbone_bd_ram_n23945, p_wishbone_bd_ram_n23946, 
        p_wishbone_bd_ram_n23947, p_wishbone_bd_ram_n23948, 
        p_wishbone_bd_ram_n23949, p_wishbone_bd_ram_n23950, 
        p_wishbone_bd_ram_n23951, p_wishbone_bd_ram_n23952, 
        p_wishbone_bd_ram_n23953, p_wishbone_bd_ram_n23954, 
        p_wishbone_bd_ram_n23955, p_wishbone_bd_ram_n23956, 
        p_wishbone_bd_ram_n23957, p_wishbone_bd_ram_n23958, 
        p_wishbone_bd_ram_n23959, p_wishbone_bd_ram_n23960, 
        p_wishbone_bd_ram_n23961, p_wishbone_bd_ram_n23962, 
        p_wishbone_bd_ram_n23963, p_wishbone_bd_ram_n23964, 
        p_wishbone_bd_ram_n23965, p_wishbone_bd_ram_n23966, 
        p_wishbone_bd_ram_n23967, p_wishbone_bd_ram_n23968, 
        p_wishbone_bd_ram_n23969, p_wishbone_bd_ram_n23970, 
        p_wishbone_bd_ram_n23971, p_wishbone_bd_ram_n23972, 
        p_wishbone_bd_ram_n23973, p_wishbone_bd_ram_n23974, 
        p_wishbone_bd_ram_n23975, p_wishbone_bd_ram_n23976, 
        p_wishbone_bd_ram_n23977, p_wishbone_bd_ram_n23978, 
        p_wishbone_bd_ram_n23979, p_wishbone_bd_ram_n23980, 
        p_wishbone_bd_ram_n23981, p_wishbone_bd_ram_n23982, 
        p_wishbone_bd_ram_n23983, p_wishbone_bd_ram_n23984, 
        p_wishbone_bd_ram_n23985, p_wishbone_bd_ram_n23986, 
        p_wishbone_bd_ram_n23987, p_wishbone_bd_ram_n23988, 
        p_wishbone_bd_ram_n23989, p_wishbone_bd_ram_n23990, 
        p_wishbone_bd_ram_n23991, p_wishbone_bd_ram_n23992, 
        p_wishbone_bd_ram_n23993, p_wishbone_bd_ram_n23994, 
        p_wishbone_bd_ram_n23995, p_wishbone_bd_ram_n23996, 
        p_wishbone_bd_ram_n23997, p_wishbone_bd_ram_n23998, 
        p_wishbone_bd_ram_n23999, p_wishbone_bd_ram_n24000, 
        p_wishbone_bd_ram_n24001, p_wishbone_bd_ram_n24002, 
        p_wishbone_bd_ram_n24003, p_wishbone_bd_ram_n24004, 
        p_wishbone_bd_ram_n24005, p_wishbone_bd_ram_n24006, 
        p_wishbone_bd_ram_n24007, p_wishbone_bd_ram_n24008, 
        p_wishbone_bd_ram_n24009, p_wishbone_bd_ram_n24010, 
        p_wishbone_bd_ram_n24011, p_wishbone_bd_ram_n24012, 
        p_wishbone_bd_ram_n24013, p_wishbone_bd_ram_n24014, 
        p_wishbone_bd_ram_n24015, p_wishbone_bd_ram_n24016, 
        p_wishbone_bd_ram_n24017, p_wishbone_bd_ram_n24018, 
        p_wishbone_bd_ram_n24019, p_wishbone_bd_ram_n24020, 
        p_wishbone_bd_ram_n24021, p_wishbone_bd_ram_n24022, 
        p_wishbone_bd_ram_n24023, p_wishbone_bd_ram_n24024, 
        p_wishbone_bd_ram_n24025, p_wishbone_bd_ram_n24026, 
        p_wishbone_bd_ram_n24027, p_wishbone_bd_ram_n24028, 
        p_wishbone_bd_ram_n24029, p_wishbone_bd_ram_n24030, 
        p_wishbone_bd_ram_n24031, p_wishbone_bd_ram_n24032, 
        p_wishbone_bd_ram_n24033, p_wishbone_bd_ram_n24034, 
        p_wishbone_bd_ram_n24035, p_wishbone_bd_ram_n24036, 
        p_wishbone_bd_ram_n24037, p_wishbone_bd_ram_n24038, 
        p_wishbone_bd_ram_n24039, p_wishbone_bd_ram_n24040, 
        p_wishbone_bd_ram_n24041, p_wishbone_bd_ram_n24042, 
        p_wishbone_bd_ram_n24043, p_wishbone_bd_ram_n24044, 
        p_wishbone_bd_ram_n24045, p_wishbone_bd_ram_n24046, 
        p_wishbone_bd_ram_n24047, p_wishbone_bd_ram_n24048, 
        p_wishbone_bd_ram_n24049, p_wishbone_bd_ram_n24050, 
        p_wishbone_bd_ram_n24051, p_wishbone_bd_ram_n24052, 
        p_wishbone_bd_ram_n24053, p_wishbone_bd_ram_n24054, 
        p_wishbone_bd_ram_n24055, p_wishbone_bd_ram_n24056, 
        p_wishbone_bd_ram_n24057, p_wishbone_bd_ram_n24058, 
        p_wishbone_bd_ram_n24059, p_wishbone_bd_ram_n24060, 
        p_wishbone_bd_ram_n24061, p_wishbone_bd_ram_n24062, 
        p_wishbone_bd_ram_n24063, p_wishbone_bd_ram_n24064, 
        p_wishbone_bd_ram_n24065, p_wishbone_bd_ram_n24066, 
        p_wishbone_bd_ram_n24067, p_wishbone_bd_ram_n24068, 
        p_wishbone_bd_ram_n24069, p_wishbone_bd_ram_n24070, 
        p_wishbone_bd_ram_n24071, p_wishbone_bd_ram_n24072, 
        p_wishbone_bd_ram_n24073, p_wishbone_bd_ram_n24074, 
        p_wishbone_bd_ram_n24075, p_wishbone_bd_ram_n24076, 
        p_wishbone_bd_ram_n24077, p_wishbone_bd_ram_n24078, 
        p_wishbone_bd_ram_n24079, p_wishbone_bd_ram_n24080, 
        p_wishbone_bd_ram_n24081, p_wishbone_bd_ram_n24082, 
        p_wishbone_bd_ram_n24083, p_wishbone_bd_ram_n24084, 
        p_wishbone_bd_ram_n24085, p_wishbone_bd_ram_n24086, 
        p_wishbone_bd_ram_n24087, p_wishbone_bd_ram_n24088, 
        p_wishbone_bd_ram_n24089, p_wishbone_bd_ram_n24090, 
        p_wishbone_bd_ram_n24091, p_wishbone_bd_ram_n24092, 
        p_wishbone_bd_ram_n24093, p_wishbone_bd_ram_n24094, 
        p_wishbone_bd_ram_n24095, p_wishbone_bd_ram_n24096, 
        p_wishbone_bd_ram_n24097, p_wishbone_bd_ram_n24098, 
        p_wishbone_bd_ram_n24099, p_wishbone_bd_ram_n24100, 
        p_wishbone_bd_ram_n24101, p_wishbone_bd_ram_n24102, 
        p_wishbone_bd_ram_n24103, p_wishbone_bd_ram_n24104, 
        p_wishbone_bd_ram_n24105, p_wishbone_bd_ram_n24106, 
        p_wishbone_bd_ram_n24107, p_wishbone_bd_ram_n24108, 
        p_wishbone_bd_ram_n24109, p_wishbone_bd_ram_n24110, 
        p_wishbone_bd_ram_n24111, p_wishbone_bd_ram_n24112, 
        p_wishbone_bd_ram_n24113, p_wishbone_bd_ram_n24114, 
        p_wishbone_bd_ram_n24115, p_wishbone_bd_ram_n24116, 
        p_wishbone_bd_ram_n24117, p_wishbone_bd_ram_n24118, 
        p_wishbone_bd_ram_n24119, p_wishbone_bd_ram_n24120, 
        p_wishbone_bd_ram_n24121, p_wishbone_bd_ram_n24122, 
        p_wishbone_bd_ram_n24123, p_wishbone_bd_ram_n24124, 
        p_wishbone_bd_ram_n24125, p_wishbone_bd_ram_n24126, 
        p_wishbone_bd_ram_n24127, p_wishbone_bd_ram_n24128, 
        p_wishbone_bd_ram_n24129, p_wishbone_bd_ram_n24130, 
        p_wishbone_bd_ram_n24131, p_wishbone_bd_ram_n24132, 
        p_wishbone_bd_ram_n24133, p_wishbone_bd_ram_n24134, 
        p_wishbone_bd_ram_n24135, p_wishbone_bd_ram_n24136, 
        p_wishbone_bd_ram_n24137, p_wishbone_bd_ram_n24138, 
        p_wishbone_bd_ram_n24139, p_wishbone_bd_ram_n24140, 
        p_wishbone_bd_ram_n24141, p_wishbone_bd_ram_n24142, 
        p_wishbone_bd_ram_n24143, p_wishbone_bd_ram_n24144, 
        p_wishbone_bd_ram_n24145, p_wishbone_bd_ram_n24146, 
        p_wishbone_bd_ram_n24147, p_wishbone_bd_ram_n24148, 
        p_wishbone_bd_ram_n24149, p_wishbone_bd_ram_n24150, 
        p_wishbone_bd_ram_n24151, p_wishbone_bd_ram_n24152, 
        p_wishbone_bd_ram_n24153, p_wishbone_bd_ram_n24154, 
        p_wishbone_bd_ram_n24155, p_wishbone_bd_ram_n24156, 
        p_wishbone_bd_ram_n24157, p_wishbone_bd_ram_n24158, 
        p_wishbone_bd_ram_n24159, p_wishbone_bd_ram_n24160, 
        p_wishbone_bd_ram_n24161, p_wishbone_bd_ram_n24162, 
        p_wishbone_bd_ram_n24163, p_wishbone_bd_ram_n24164, 
        p_wishbone_bd_ram_n24165, p_wishbone_bd_ram_n24166, 
        p_wishbone_bd_ram_n24167, p_wishbone_bd_ram_n24168, 
        p_wishbone_bd_ram_n24169, p_wishbone_bd_ram_n24170, 
        p_wishbone_bd_ram_n24171, p_wishbone_bd_ram_n24172, 
        p_wishbone_bd_ram_n24173, p_wishbone_bd_ram_n24174, 
        p_wishbone_bd_ram_n24175, p_wishbone_bd_ram_n24176, 
        p_wishbone_bd_ram_n24177, p_wishbone_bd_ram_n24178, 
        p_wishbone_bd_ram_n24179, p_wishbone_bd_ram_n24180, 
        p_wishbone_bd_ram_n24181, p_wishbone_bd_ram_n24182, 
        p_wishbone_bd_ram_n24183, p_wishbone_bd_ram_n24184, 
        p_wishbone_bd_ram_n24185, p_wishbone_bd_ram_n24186, 
        p_wishbone_bd_ram_n24187, p_wishbone_bd_ram_n24188, 
        p_wishbone_bd_ram_n24189, p_wishbone_bd_ram_n24190, 
        p_wishbone_bd_ram_n24191, p_wishbone_bd_ram_n24192, 
        p_wishbone_bd_ram_n24193, p_wishbone_bd_ram_n24194, 
        p_wishbone_bd_ram_n24195, p_wishbone_bd_ram_n24196, 
        p_wishbone_bd_ram_n24197, p_wishbone_bd_ram_n24198, 
        p_wishbone_bd_ram_n24199, p_wishbone_bd_ram_n24200, 
        p_wishbone_bd_ram_n24201, p_wishbone_bd_ram_n24202, 
        p_wishbone_bd_ram_n24203, p_wishbone_bd_ram_n24204, 
        p_wishbone_bd_ram_n24205, p_wishbone_bd_ram_n24206, 
        p_wishbone_bd_ram_n24207, p_wishbone_bd_ram_n24208, 
        p_wishbone_bd_ram_n24209, p_wishbone_bd_ram_n24210, 
        p_wishbone_bd_ram_n24211, p_wishbone_bd_ram_n24212, 
        p_wishbone_bd_ram_n24213, p_wishbone_bd_ram_n24214, 
        p_wishbone_bd_ram_n24215, p_wishbone_bd_ram_n24216, 
        p_wishbone_bd_ram_n24217, p_wishbone_bd_ram_n24218, 
        p_wishbone_bd_ram_n24219, p_wishbone_bd_ram_n24220, 
        p_wishbone_bd_ram_n24221, p_wishbone_bd_ram_n24222, 
        p_wishbone_bd_ram_n24223, p_wishbone_bd_ram_n24224, 
        p_wishbone_bd_ram_n24225, p_wishbone_bd_ram_n24226, 
        p_wishbone_bd_ram_n24227, p_wishbone_bd_ram_n24228, 
        p_wishbone_bd_ram_n24229, p_wishbone_bd_ram_n24230, 
        p_wishbone_bd_ram_n24231, p_wishbone_bd_ram_n24232, 
        p_wishbone_bd_ram_n24233, p_wishbone_bd_ram_n24234, 
        p_wishbone_bd_ram_n24235, p_wishbone_bd_ram_n24236, 
        p_wishbone_bd_ram_n24237, p_wishbone_bd_ram_n24238, 
        p_wishbone_bd_ram_n24239, p_wishbone_bd_ram_n24240, 
        p_wishbone_bd_ram_n24241, p_wishbone_bd_ram_n24242, 
        p_wishbone_bd_ram_n24243, p_wishbone_bd_ram_n24244, 
        p_wishbone_bd_ram_n24245, p_wishbone_bd_ram_n24246, 
        p_wishbone_bd_ram_n24247, p_wishbone_bd_ram_n24248, 
        p_wishbone_bd_ram_n24249, p_wishbone_bd_ram_n24250, 
        p_wishbone_bd_ram_n24251, p_wishbone_bd_ram_n24252, 
        p_wishbone_bd_ram_n24253, p_wishbone_bd_ram_n24254, 
        p_wishbone_bd_ram_n24255, p_wishbone_bd_ram_n24256, 
        p_wishbone_bd_ram_n24257, p_wishbone_bd_ram_n24258, 
        p_wishbone_bd_ram_n24259, p_wishbone_bd_ram_n24260, 
        p_wishbone_bd_ram_n24261, p_wishbone_bd_ram_n24262, 
        p_wishbone_bd_ram_n24263, p_wishbone_bd_ram_n24264, 
        p_wishbone_bd_ram_n24265, p_wishbone_bd_ram_n24266, 
        p_wishbone_bd_ram_n24267, p_wishbone_bd_ram_n24268, 
        p_wishbone_bd_ram_n24269, p_wishbone_bd_ram_n24270, 
        p_wishbone_bd_ram_n24271, p_wishbone_bd_ram_n24272, 
        p_wishbone_bd_ram_n24273, p_wishbone_bd_ram_n24274, 
        p_wishbone_bd_ram_n24275, p_wishbone_bd_ram_n24276, 
        p_wishbone_bd_ram_n24277, p_wishbone_bd_ram_n24278, 
        p_wishbone_bd_ram_n24279, p_wishbone_bd_ram_n24280, 
        p_wishbone_bd_ram_n24281, p_wishbone_bd_ram_n24282, 
        p_wishbone_bd_ram_n24283, p_wishbone_bd_ram_n24284, 
        p_wishbone_bd_ram_n24285, p_wishbone_bd_ram_n24286, 
        p_wishbone_bd_ram_n24287, p_wishbone_bd_ram_n24288, 
        p_wishbone_bd_ram_n24289, p_wishbone_bd_ram_n24290, 
        p_wishbone_bd_ram_n24291, p_wishbone_bd_ram_n24292, 
        p_wishbone_bd_ram_n24293, p_wishbone_bd_ram_n24294, 
        p_wishbone_bd_ram_n24295, p_wishbone_bd_ram_n24296, 
        p_wishbone_bd_ram_n24297, p_wishbone_bd_ram_n24298, 
        p_wishbone_bd_ram_n24299, p_wishbone_bd_ram_n24300, 
        p_wishbone_bd_ram_n24301, p_wishbone_bd_ram_n24302, 
        p_wishbone_bd_ram_n24303, p_wishbone_bd_ram_n24304, 
        p_wishbone_bd_ram_n24305, p_wishbone_bd_ram_n24306, 
        p_wishbone_bd_ram_n24307, p_wishbone_bd_ram_n24308, 
        p_wishbone_bd_ram_n24309, p_wishbone_bd_ram_n24310, 
        p_wishbone_bd_ram_n24311, p_wishbone_bd_ram_n24312, 
        p_wishbone_bd_ram_n24313, p_wishbone_bd_ram_n24314, 
        p_wishbone_bd_ram_n24315, p_wishbone_bd_ram_n24316, 
        p_wishbone_bd_ram_n24317, p_wishbone_bd_ram_n24318, 
        p_wishbone_bd_ram_n24319, p_wishbone_bd_ram_n24320, 
        p_wishbone_bd_ram_n24321, p_wishbone_bd_ram_n24322, 
        p_wishbone_bd_ram_n24323, p_wishbone_bd_ram_n24324, 
        p_wishbone_bd_ram_n24325, p_wishbone_bd_ram_n24326, 
        p_wishbone_bd_ram_n24327, p_wishbone_bd_ram_n24328, 
        p_wishbone_bd_ram_n24329, p_wishbone_bd_ram_n24330, 
        p_wishbone_bd_ram_n24331, p_wishbone_bd_ram_n24332, 
        p_wishbone_bd_ram_n24333, p_wishbone_bd_ram_n24334, 
        p_wishbone_bd_ram_n24335, p_wishbone_bd_ram_n24336, 
        p_wishbone_bd_ram_n24337, p_wishbone_bd_ram_n24338, 
        p_wishbone_bd_ram_n24339, p_wishbone_bd_ram_n24340, 
        p_wishbone_bd_ram_n24341, p_wishbone_bd_ram_n24342, 
        p_wishbone_bd_ram_n24343, p_wishbone_bd_ram_n24344, 
        p_wishbone_bd_ram_n24345, p_wishbone_bd_ram_n24346, 
        p_wishbone_bd_ram_n24347, p_wishbone_bd_ram_n24348, 
        p_wishbone_bd_ram_n24349, p_wishbone_bd_ram_n24350, 
        p_wishbone_bd_ram_n24351, p_wishbone_bd_ram_n24352, 
        p_wishbone_bd_ram_n24353, p_wishbone_bd_ram_n24354, 
        p_wishbone_bd_ram_n24355, p_wishbone_bd_ram_n24356, 
        p_wishbone_bd_ram_n24357, p_wishbone_bd_ram_n24358, 
        p_wishbone_bd_ram_n24359, p_wishbone_bd_ram_n24360, 
        p_wishbone_bd_ram_n24361, p_wishbone_bd_ram_n24362, 
        p_wishbone_bd_ram_n24363, p_wishbone_bd_ram_n24364, 
        p_wishbone_bd_ram_n24365, p_wishbone_bd_ram_n24366, 
        p_wishbone_bd_ram_n24367, p_wishbone_bd_ram_n24368, 
        p_wishbone_bd_ram_n24369, p_wishbone_bd_ram_n24370, 
        p_wishbone_bd_ram_n24371, p_wishbone_bd_ram_n24372, 
        p_wishbone_bd_ram_n24373, p_wishbone_bd_ram_n24374, 
        p_wishbone_bd_ram_n24375, p_wishbone_bd_ram_n24376, 
        p_wishbone_bd_ram_n24377, p_wishbone_bd_ram_n24378, 
        p_wishbone_bd_ram_n24379, p_wishbone_bd_ram_n24380, 
        p_wishbone_bd_ram_n24381, p_wishbone_bd_ram_n24382, 
        p_wishbone_bd_ram_n24383, p_wishbone_bd_ram_n24384, 
        p_wishbone_bd_ram_n24385, p_wishbone_bd_ram_n24386, 
        p_wishbone_bd_ram_n24387, p_wishbone_bd_ram_n24388, 
        p_wishbone_bd_ram_n24389, p_wishbone_bd_ram_n24390, 
        p_wishbone_bd_ram_n24391, p_wishbone_bd_ram_n24392, 
        p_wishbone_bd_ram_n24393, p_wishbone_bd_ram_n24394, 
        p_wishbone_bd_ram_n24395, p_wishbone_bd_ram_n24396, 
        p_wishbone_bd_ram_n24397, p_wishbone_bd_ram_n24398, 
        p_wishbone_bd_ram_n24399, p_wishbone_bd_ram_n24400, 
        p_wishbone_bd_ram_n24401, p_wishbone_bd_ram_n24402, 
        p_wishbone_bd_ram_n24403, p_wishbone_bd_ram_n24404, 
        p_wishbone_bd_ram_n24405, p_wishbone_bd_ram_n24406, 
        p_wishbone_bd_ram_n24407, p_wishbone_bd_ram_n24408, 
        p_wishbone_bd_ram_n24409, p_wishbone_bd_ram_n24410, 
        p_wishbone_bd_ram_n24411, p_wishbone_bd_ram_n24412, 
        p_wishbone_bd_ram_n24413, p_wishbone_bd_ram_n24414, 
        p_wishbone_bd_ram_n24415, p_wishbone_bd_ram_n24416, 
        p_wishbone_bd_ram_n24417, p_wishbone_bd_ram_n24418, 
        p_wishbone_bd_ram_n24419, p_wishbone_bd_ram_n24420, 
        p_wishbone_bd_ram_n24421, p_wishbone_bd_ram_n24422, 
        p_wishbone_bd_ram_n24423, p_wishbone_bd_ram_n24424, 
        p_wishbone_bd_ram_n24425, p_wishbone_bd_ram_n24426, 
        p_wishbone_bd_ram_n24427, p_wishbone_bd_ram_n24428, 
        p_wishbone_bd_ram_n24429, p_wishbone_bd_ram_n24430, 
        p_wishbone_bd_ram_n24431, p_wishbone_bd_ram_n24432, 
        p_wishbone_bd_ram_n24433, p_wishbone_bd_ram_n24434, 
        p_wishbone_bd_ram_n24435, p_wishbone_bd_ram_n24436, 
        p_wishbone_bd_ram_n24437, p_wishbone_bd_ram_n24438, 
        p_wishbone_bd_ram_n24439, p_wishbone_bd_ram_n24440, 
        p_wishbone_bd_ram_n24441, p_wishbone_bd_ram_n24442, 
        p_wishbone_bd_ram_n24443, p_wishbone_bd_ram_n24444, 
        p_wishbone_bd_ram_n24445, p_wishbone_bd_ram_n24446, 
        p_wishbone_bd_ram_n24447, p_wishbone_bd_ram_n24448, 
        p_wishbone_bd_ram_n24449, p_wishbone_bd_ram_n24450, 
        p_wishbone_bd_ram_n24451, p_wishbone_bd_ram_n24452, 
        p_wishbone_bd_ram_n24453, p_wishbone_bd_ram_n24454, 
        p_wishbone_bd_ram_n24455, p_wishbone_bd_ram_n24456, 
        p_wishbone_bd_ram_n24457, p_wishbone_bd_ram_n24458, 
        p_wishbone_bd_ram_n24459, p_wishbone_bd_ram_n24460, 
        p_wishbone_bd_ram_n24461, p_wishbone_bd_ram_n24462, 
        p_wishbone_bd_ram_n24463, p_wishbone_bd_ram_n24464, 
        p_wishbone_bd_ram_n24465, p_wishbone_bd_ram_n24466, 
        p_wishbone_bd_ram_n24467, p_wishbone_bd_ram_n24468, 
        p_wishbone_bd_ram_n24469, p_wishbone_bd_ram_n24470, 
        p_wishbone_bd_ram_n24471, p_wishbone_bd_ram_n24472, 
        p_wishbone_bd_ram_n24473, p_wishbone_bd_ram_n24474, 
        p_wishbone_bd_ram_n24475, p_wishbone_bd_ram_n24476, 
        p_wishbone_bd_ram_n24477, p_wishbone_bd_ram_n24478, 
        p_wishbone_bd_ram_n24479, p_wishbone_bd_ram_n24480, 
        p_wishbone_bd_ram_n24481, p_wishbone_bd_ram_n24482, 
        p_wishbone_bd_ram_n24483, p_wishbone_bd_ram_n24484, 
        p_wishbone_bd_ram_n24485, p_wishbone_bd_ram_n24486, 
        p_wishbone_bd_ram_n24487, p_wishbone_bd_ram_n24488, 
        p_wishbone_bd_ram_n24489, p_wishbone_bd_ram_n24490, 
        p_wishbone_bd_ram_n24491, p_wishbone_bd_ram_n24492, 
        p_wishbone_bd_ram_n24493, p_wishbone_bd_ram_n24494, 
        p_wishbone_bd_ram_n24495, p_wishbone_bd_ram_n24496, 
        p_wishbone_bd_ram_n24497, p_wishbone_bd_ram_n24498, 
        p_wishbone_bd_ram_n24499, p_wishbone_bd_ram_n24500, 
        p_wishbone_bd_ram_n24501, p_wishbone_bd_ram_n24502, 
        p_wishbone_bd_ram_n24503, p_wishbone_bd_ram_n24504, 
        p_wishbone_bd_ram_n24505, p_wishbone_bd_ram_n24506, 
        p_wishbone_bd_ram_n24507, p_wishbone_bd_ram_n24508, 
        p_wishbone_bd_ram_n24509, p_wishbone_bd_ram_n24510, 
        p_wishbone_bd_ram_n24511, p_wishbone_bd_ram_n24512, 
        p_wishbone_bd_ram_n24513, p_wishbone_bd_ram_n24514, 
        p_wishbone_bd_ram_n24515, p_wishbone_bd_ram_n24516, 
        p_wishbone_bd_ram_n24517, p_wishbone_bd_ram_n24518, 
        p_wishbone_bd_ram_n24519, p_wishbone_bd_ram_n24520, 
        p_wishbone_bd_ram_n24521, p_wishbone_bd_ram_n24522, 
        p_wishbone_bd_ram_n24523, p_wishbone_bd_ram_n24524, 
        p_wishbone_bd_ram_n24525, p_wishbone_bd_ram_n24526, 
        p_wishbone_bd_ram_n24527, p_wishbone_bd_ram_n24528, 
        p_wishbone_bd_ram_n24529, p_wishbone_bd_ram_n24530, 
        p_wishbone_bd_ram_n24531, p_wishbone_bd_ram_n24532, 
        p_wishbone_bd_ram_n24533, p_wishbone_bd_ram_n24534, 
        p_wishbone_bd_ram_n24535, p_wishbone_bd_ram_n24536, 
        p_wishbone_bd_ram_n24537, p_wishbone_bd_ram_n24538, 
        p_wishbone_bd_ram_n24539, p_wishbone_bd_ram_n24540, 
        p_wishbone_bd_ram_n24541, p_wishbone_bd_ram_n24542, 
        p_wishbone_bd_ram_n24543, p_wishbone_bd_ram_n24544, 
        p_wishbone_bd_ram_n24545, p_wishbone_bd_ram_n24546, 
        p_wishbone_bd_ram_n24547, p_wishbone_bd_ram_n24548, 
        p_wishbone_bd_ram_n24549, p_wishbone_bd_ram_n24550, 
        p_wishbone_bd_ram_n24551, p_wishbone_bd_ram_n24552, 
        p_wishbone_bd_ram_n24553, p_wishbone_bd_ram_n24554, 
        p_wishbone_bd_ram_n24555, p_wishbone_bd_ram_n24556, 
        p_wishbone_bd_ram_n24557, p_wishbone_bd_ram_n24558, 
        p_wishbone_bd_ram_n24559, p_wishbone_bd_ram_n24560, 
        p_wishbone_bd_ram_n24561, p_wishbone_bd_ram_n24562, 
        p_wishbone_bd_ram_n24563, p_wishbone_bd_ram_n24564, 
        p_wishbone_bd_ram_n24565, p_wishbone_bd_ram_n24566, 
        p_wishbone_bd_ram_n24567, p_wishbone_bd_ram_n24568, 
        p_wishbone_bd_ram_n24569, p_wishbone_bd_ram_n24570, 
        p_wishbone_bd_ram_n24571, p_wishbone_bd_ram_n24572, 
        p_wishbone_bd_ram_n24573, p_wishbone_bd_ram_n24574, 
        p_wishbone_bd_ram_n24575, p_wishbone_bd_ram_n24576, 
        p_wishbone_bd_ram_n24577, p_wishbone_bd_ram_n24578, 
        p_wishbone_bd_ram_n24579, p_wishbone_bd_ram_n24580, 
        p_wishbone_bd_ram_n24581, p_wishbone_bd_ram_n24582, 
        p_wishbone_bd_ram_n24583, p_wishbone_bd_ram_n24584, 
        p_wishbone_bd_ram_n24585, p_wishbone_bd_ram_n24586, 
        p_wishbone_bd_ram_n24587, p_wishbone_bd_ram_n24588, 
        p_wishbone_bd_ram_n24589, p_wishbone_bd_ram_n24590, 
        p_wishbone_bd_ram_n24591, p_wishbone_bd_ram_n24592, 
        p_wishbone_bd_ram_n24593, p_wishbone_bd_ram_n24594, 
        p_wishbone_bd_ram_n24595, p_wishbone_bd_ram_n24596, 
        p_wishbone_bd_ram_n24597, p_wishbone_bd_ram_n24598, 
        p_wishbone_bd_ram_n24599, p_wishbone_bd_ram_n24600, 
        p_wishbone_bd_ram_n24601, p_wishbone_bd_ram_n24602, 
        p_wishbone_bd_ram_n24603, p_wishbone_bd_ram_n24604, 
        p_wishbone_bd_ram_n24605, p_wishbone_bd_ram_n24606, 
        p_wishbone_bd_ram_n24607, p_wishbone_bd_ram_n24608, 
        p_wishbone_bd_ram_n24609, p_wishbone_bd_ram_n24610, 
        p_wishbone_bd_ram_n24611, p_wishbone_bd_ram_n24612, 
        p_wishbone_bd_ram_n24613, p_wishbone_bd_ram_n24614, 
        p_wishbone_bd_ram_n24615, p_wishbone_bd_ram_n24616, 
        p_wishbone_bd_ram_n24617, p_wishbone_bd_ram_n24618, 
        p_wishbone_bd_ram_n24619, p_wishbone_bd_ram_n24620, 
        p_wishbone_bd_ram_n24621, p_wishbone_bd_ram_n24622, 
        p_wishbone_bd_ram_n24623, p_wishbone_bd_ram_n24624, 
        p_wishbone_bd_ram_n24625, p_wishbone_bd_ram_n24626, 
        p_wishbone_bd_ram_n24627, p_wishbone_bd_ram_n24628, 
        p_wishbone_bd_ram_n24629, p_wishbone_bd_ram_n24630, 
        p_wishbone_bd_ram_n24631, p_wishbone_bd_ram_n24632, 
        p_wishbone_bd_ram_n24633, p_wishbone_bd_ram_n24634, 
        p_wishbone_bd_ram_n24635, p_wishbone_bd_ram_n24636, 
        p_wishbone_bd_ram_n24637, p_wishbone_bd_ram_n24638, 
        p_wishbone_bd_ram_n24639, p_wishbone_bd_ram_n24640, 
        p_wishbone_bd_ram_n24641, p_wishbone_bd_ram_n24642, 
        p_wishbone_bd_ram_n24643, p_wishbone_bd_ram_n24644, 
        p_wishbone_bd_ram_n24645, p_wishbone_bd_ram_n24646, 
        p_wishbone_bd_ram_n24647, p_wishbone_bd_ram_n24648, 
        p_wishbone_bd_ram_n24649, p_wishbone_bd_ram_n24650, 
        p_wishbone_bd_ram_n24651, p_wishbone_bd_ram_n24652, 
        p_wishbone_bd_ram_n24653, p_wishbone_bd_ram_n24654, 
        p_wishbone_bd_ram_n24655, p_wishbone_bd_ram_n24656, 
        p_wishbone_bd_ram_n24657, p_wishbone_bd_ram_n24658, 
        p_wishbone_bd_ram_n24659, p_wishbone_bd_ram_n24660, 
        p_wishbone_bd_ram_n24661, p_wishbone_bd_ram_n24662, 
        p_wishbone_bd_ram_n24663, p_wishbone_bd_ram_n24664, 
        p_wishbone_bd_ram_n24665, p_wishbone_bd_ram_n24666, 
        p_wishbone_bd_ram_n24667, p_wishbone_bd_ram_n24668, 
        p_wishbone_bd_ram_n24669, p_wishbone_bd_ram_n24670, 
        p_wishbone_bd_ram_n24671, p_wishbone_bd_ram_n24672, 
        p_wishbone_bd_ram_n24673, p_wishbone_bd_ram_n24674, 
        p_wishbone_bd_ram_n24675, p_wishbone_bd_ram_n24676, 
        p_wishbone_bd_ram_n24677, p_wishbone_bd_ram_n24678, 
        p_wishbone_bd_ram_n24679, p_wishbone_bd_ram_n24680, 
        p_wishbone_bd_ram_n24681, p_wishbone_bd_ram_n24682, 
        p_wishbone_bd_ram_n24683, p_wishbone_bd_ram_n24684, 
        p_wishbone_bd_ram_n24685, p_wishbone_bd_ram_n24686, 
        p_wishbone_bd_ram_n24687, p_wishbone_bd_ram_n24688, 
        p_wishbone_bd_ram_n24689, p_wishbone_bd_ram_n24690, 
        p_wishbone_bd_ram_n24691, p_wishbone_bd_ram_n24692, 
        p_wishbone_bd_ram_n24693, p_wishbone_bd_ram_n24694, 
        p_wishbone_bd_ram_n24695, p_wishbone_bd_ram_n24696, 
        p_wishbone_bd_ram_n24697, p_wishbone_bd_ram_n24698, 
        p_wishbone_bd_ram_n24699, p_wishbone_bd_ram_n24700, 
        p_wishbone_bd_ram_n24701, p_wishbone_bd_ram_n24702, 
        p_wishbone_bd_ram_n24703, p_wishbone_bd_ram_n24704, 
        p_wishbone_bd_ram_n24705, p_wishbone_bd_ram_n24706, 
        p_wishbone_bd_ram_n24707, p_wishbone_bd_ram_n24708, 
        p_wishbone_bd_ram_n24709, p_wishbone_bd_ram_n24710, 
        p_wishbone_bd_ram_n24711, p_wishbone_bd_ram_n24712, 
        p_wishbone_bd_ram_n24713, p_wishbone_bd_ram_n24714, 
        p_wishbone_bd_ram_n24715, p_wishbone_bd_ram_n24716, 
        p_wishbone_bd_ram_n24717, p_wishbone_bd_ram_n24718, 
        p_wishbone_bd_ram_n24719, p_wishbone_bd_ram_n24720, 
        p_wishbone_bd_ram_n24721, p_wishbone_bd_ram_n24722, 
        p_wishbone_bd_ram_n24723, p_wishbone_bd_ram_n24724, 
        p_wishbone_bd_ram_n24725, p_wishbone_bd_ram_n24726, 
        p_wishbone_bd_ram_n24727, p_wishbone_bd_ram_n24728, 
        p_wishbone_bd_ram_n24729, p_wishbone_bd_ram_n24730, 
        p_wishbone_bd_ram_n24731, p_wishbone_bd_ram_n24732, 
        p_wishbone_bd_ram_n24733, p_wishbone_bd_ram_n24734, 
        p_wishbone_bd_ram_n24735, p_wishbone_bd_ram_n24736, 
        p_wishbone_bd_ram_n24737, p_wishbone_bd_ram_n24738, 
        p_wishbone_bd_ram_n24739, p_wishbone_bd_ram_n24740, 
        p_wishbone_bd_ram_n24741, p_wishbone_bd_ram_n24742, 
        p_wishbone_bd_ram_n24743, p_wishbone_bd_ram_n24744, 
        p_wishbone_bd_ram_n24745, p_wishbone_bd_ram_n24746, 
        p_wishbone_bd_ram_n24747, p_wishbone_bd_ram_n24748, 
        p_wishbone_bd_ram_n24749, p_wishbone_bd_ram_n24750, 
        p_wishbone_bd_ram_n24751, p_wishbone_bd_ram_n24752, 
        p_wishbone_bd_ram_n24753, p_wishbone_bd_ram_n24754, 
        p_wishbone_bd_ram_n24755, p_wishbone_bd_ram_n24756, 
        p_wishbone_bd_ram_n24757, p_wishbone_bd_ram_n24758, 
        p_wishbone_bd_ram_n24759, p_wishbone_bd_ram_n24760, 
        p_wishbone_bd_ram_n24761, p_wishbone_bd_ram_n24762, 
        p_wishbone_bd_ram_n24763, p_wishbone_bd_ram_n24764, 
        p_wishbone_bd_ram_n24765, p_wishbone_bd_ram_n24766, 
        p_wishbone_bd_ram_n24767, p_wishbone_bd_ram_n24768, 
        p_wishbone_bd_ram_n24769, p_wishbone_bd_ram_n24770, 
        p_wishbone_bd_ram_n24771, p_wishbone_bd_ram_n24772, 
        p_wishbone_bd_ram_n24773, p_wishbone_bd_ram_n24774, 
        p_wishbone_bd_ram_n24775, p_wishbone_bd_ram_n24776, 
        p_wishbone_bd_ram_n24777, p_wishbone_bd_ram_n24778, 
        p_wishbone_bd_ram_n24779, p_wishbone_bd_ram_n24780, 
        p_wishbone_bd_ram_n24781, p_wishbone_bd_ram_n24782, 
        p_wishbone_bd_ram_n24783, p_wishbone_bd_ram_n24784, 
        p_wishbone_bd_ram_n24785, p_wishbone_bd_ram_n24786, 
        p_wishbone_bd_ram_n24787, p_wishbone_bd_ram_n24788, 
        p_wishbone_bd_ram_n24789, p_wishbone_bd_ram_n24790, 
        p_wishbone_bd_ram_n24791, p_wishbone_bd_ram_n24792, 
        p_wishbone_bd_ram_n24793, p_wishbone_bd_ram_n24794, 
        p_wishbone_bd_ram_n24795, p_wishbone_bd_ram_n24796, 
        p_wishbone_bd_ram_n24797, p_wishbone_bd_ram_n24798, 
        p_wishbone_bd_ram_n24799, p_wishbone_bd_ram_n24800, 
        p_wishbone_bd_ram_n24801, p_wishbone_bd_ram_n24802, 
        p_wishbone_bd_ram_n24803, p_wishbone_bd_ram_n24804, 
        p_wishbone_bd_ram_n24805, p_wishbone_bd_ram_n24806, 
        p_wishbone_bd_ram_n24807, p_wishbone_bd_ram_n24808, 
        p_wishbone_bd_ram_n24809, p_wishbone_bd_ram_n24810, 
        p_wishbone_bd_ram_n24811, p_wishbone_bd_ram_n24812, 
        p_wishbone_bd_ram_n24813, p_wishbone_bd_ram_n24814, 
        p_wishbone_bd_ram_n24815, p_wishbone_bd_ram_n24816, 
        p_wishbone_bd_ram_n24817, p_wishbone_bd_ram_n24818, 
        p_wishbone_bd_ram_n24819, p_wishbone_bd_ram_n24820, 
        p_wishbone_bd_ram_n24821, p_wishbone_bd_ram_n24822, 
        p_wishbone_bd_ram_n24823, p_wishbone_bd_ram_n24824, 
        p_wishbone_bd_ram_n24825, p_wishbone_bd_ram_n24826, 
        p_wishbone_bd_ram_n24827, p_wishbone_bd_ram_n24828, 
        p_wishbone_bd_ram_n24829, p_wishbone_bd_ram_n24830, 
        p_wishbone_bd_ram_n24831, p_wishbone_bd_ram_n24832, 
        p_wishbone_bd_ram_n24833, p_wishbone_bd_ram_n24834, 
        p_wishbone_bd_ram_n24835, p_wishbone_bd_ram_n24836, 
        p_wishbone_bd_ram_n24837, p_wishbone_bd_ram_n24838, 
        p_wishbone_bd_ram_n24839, p_wishbone_bd_ram_n24840, 
        p_wishbone_bd_ram_n24841, p_wishbone_bd_ram_n24842, 
        p_wishbone_bd_ram_n24843, p_wishbone_bd_ram_n24844, 
        p_wishbone_bd_ram_n24845, p_wishbone_bd_ram_n24846, 
        p_wishbone_bd_ram_n24847, p_wishbone_bd_ram_n24848, 
        p_wishbone_bd_ram_n24849, p_wishbone_bd_ram_n24850, 
        p_wishbone_bd_ram_n24851, p_wishbone_bd_ram_n24852, 
        p_wishbone_bd_ram_n24853, p_wishbone_bd_ram_n24854, 
        p_wishbone_bd_ram_n24855, p_wishbone_bd_ram_n24856, 
        p_wishbone_bd_ram_n24857, p_wishbone_bd_ram_n24858, 
        p_wishbone_bd_ram_n24859, p_wishbone_bd_ram_n24860, 
        p_wishbone_bd_ram_n24861, p_wishbone_bd_ram_n24862, 
        p_wishbone_bd_ram_n24863, p_wishbone_bd_ram_n24864, 
        p_wishbone_bd_ram_n24865, p_wishbone_bd_ram_n24866, 
        p_wishbone_bd_ram_n24867, p_wishbone_bd_ram_n24868, 
        p_wishbone_bd_ram_n24869, p_wishbone_bd_ram_n24870, 
        p_wishbone_bd_ram_n24871, p_wishbone_bd_ram_n24872, 
        p_wishbone_bd_ram_n24873, p_wishbone_bd_ram_n24874, 
        p_wishbone_bd_ram_n24875, p_wishbone_bd_ram_n24876, 
        p_wishbone_bd_ram_n24877, p_wishbone_bd_ram_n24878, 
        p_wishbone_bd_ram_n24879, p_wishbone_bd_ram_n24880, 
        p_wishbone_bd_ram_n24881, p_wishbone_bd_ram_n24882, 
        p_wishbone_bd_ram_n24883, p_wishbone_bd_ram_n24884, 
        p_wishbone_bd_ram_n24885, p_wishbone_bd_ram_n24886, 
        p_wishbone_bd_ram_n24887, p_wishbone_bd_ram_n24888, 
        p_wishbone_bd_ram_n24889, p_wishbone_bd_ram_n24890, 
        p_wishbone_bd_ram_n24891, p_wishbone_bd_ram_n24892, 
        p_wishbone_bd_ram_n24893, p_wishbone_bd_ram_n24894, 
        p_wishbone_bd_ram_n24895, p_wishbone_bd_ram_n24896, 
        p_wishbone_bd_ram_n24897, p_wishbone_bd_ram_n24898, 
        p_wishbone_bd_ram_n24899, p_wishbone_bd_ram_n24900, 
        p_wishbone_bd_ram_n24901, p_wishbone_bd_ram_n24902, 
        p_wishbone_bd_ram_n24903, p_wishbone_bd_ram_n24904, 
        p_wishbone_bd_ram_n24905, p_wishbone_bd_ram_n24906, 
        p_wishbone_bd_ram_n24907, p_wishbone_bd_ram_n24908, 
        p_wishbone_bd_ram_n24909, p_wishbone_bd_ram_n24910, 
        p_wishbone_bd_ram_n24911, p_wishbone_bd_ram_n24912, 
        p_wishbone_bd_ram_n24913, p_wishbone_bd_ram_n24914, 
        p_wishbone_bd_ram_n24915, p_wishbone_bd_ram_n24916, 
        p_wishbone_bd_ram_n24917, p_wishbone_bd_ram_n24918, 
        p_wishbone_bd_ram_n24919, p_wishbone_bd_ram_n24920, 
        p_wishbone_bd_ram_n24921, p_wishbone_bd_ram_n24922, 
        p_wishbone_bd_ram_n24923, p_wishbone_bd_ram_n24924, 
        p_wishbone_bd_ram_n24925, p_wishbone_bd_ram_n24926, 
        p_wishbone_bd_ram_n24927, p_wishbone_bd_ram_n24928, 
        p_wishbone_bd_ram_n24929, p_wishbone_bd_ram_n24930, 
        p_wishbone_bd_ram_n24931, p_wishbone_bd_ram_n24932, 
        p_wishbone_bd_ram_n24933, p_wishbone_bd_ram_n24934, 
        p_wishbone_bd_ram_n24935, p_wishbone_bd_ram_n24936, 
        p_wishbone_bd_ram_n24937, p_wishbone_bd_ram_n24938, 
        p_wishbone_bd_ram_n24939, p_wishbone_bd_ram_n24940, 
        p_wishbone_bd_ram_n24941, p_wishbone_bd_ram_n24942, 
        p_wishbone_bd_ram_n24943, p_wishbone_bd_ram_n24944, 
        p_wishbone_bd_ram_n24945, p_wishbone_bd_ram_n24946, 
        p_wishbone_bd_ram_n24947, p_wishbone_bd_ram_n24948, 
        p_wishbone_bd_ram_n24949, p_wishbone_bd_ram_n24950, 
        p_wishbone_bd_ram_n24951, p_wishbone_bd_ram_n24952, 
        p_wishbone_bd_ram_n24953, p_wishbone_bd_ram_n24954, 
        p_wishbone_bd_ram_n24955, p_wishbone_bd_ram_n24956, 
        p_wishbone_bd_ram_n24957, p_wishbone_bd_ram_n24958, 
        p_wishbone_bd_ram_n24959, p_wishbone_bd_ram_n24960, 
        p_wishbone_bd_ram_n24961, p_wishbone_bd_ram_n24962, 
        p_wishbone_bd_ram_n24963, p_wishbone_bd_ram_n24964, 
        p_wishbone_bd_ram_n24965, p_wishbone_bd_ram_n24966, 
        p_wishbone_bd_ram_n24967, p_wishbone_bd_ram_n24968, 
        p_wishbone_bd_ram_n24969, p_wishbone_bd_ram_n24970, 
        p_wishbone_bd_ram_n24971, p_wishbone_bd_ram_n24972, 
        p_wishbone_bd_ram_n24973, p_wishbone_bd_ram_n24974, 
        p_wishbone_bd_ram_n24975, p_wishbone_bd_ram_n24976, 
        p_wishbone_bd_ram_n24977, p_wishbone_bd_ram_n24978, 
        p_wishbone_bd_ram_n24979, p_wishbone_bd_ram_n24980, 
        p_wishbone_bd_ram_n24981, p_wishbone_bd_ram_n24982, 
        p_wishbone_bd_ram_n24983, p_wishbone_bd_ram_n24984, 
        p_wishbone_bd_ram_n24985, p_wishbone_bd_ram_n24986, 
        p_wishbone_bd_ram_n24987, p_wishbone_bd_ram_n24988, 
        p_wishbone_bd_ram_n24989, p_wishbone_bd_ram_n24990, 
        p_wishbone_bd_ram_n24991, p_wishbone_bd_ram_n24992, 
        p_wishbone_bd_ram_n24993, p_wishbone_bd_ram_n24994, 
        p_wishbone_bd_ram_n24995, p_wishbone_bd_ram_n24996, 
        p_wishbone_bd_ram_n24997, p_wishbone_bd_ram_n24998, 
        p_wishbone_bd_ram_n24999, p_wishbone_bd_ram_n25000, 
        p_wishbone_bd_ram_n25001, p_wishbone_bd_ram_n25002, 
        p_wishbone_bd_ram_n25003, p_wishbone_bd_ram_n25004, 
        p_wishbone_bd_ram_n25005, p_wishbone_bd_ram_n25006, 
        p_wishbone_bd_ram_n25007, p_wishbone_bd_ram_n25008, 
        p_wishbone_bd_ram_n25009, p_wishbone_bd_ram_n25010, 
        p_wishbone_bd_ram_n25011, p_wishbone_bd_ram_n25012, 
        p_wishbone_bd_ram_n25013, p_wishbone_bd_ram_n25014, 
        p_wishbone_bd_ram_n25015, p_wishbone_bd_ram_n25016, 
        p_wishbone_bd_ram_n25017, p_wishbone_bd_ram_n25018, 
        p_wishbone_bd_ram_n25019, p_wishbone_bd_ram_n25020, 
        p_wishbone_bd_ram_n25021, p_wishbone_bd_ram_n25022, 
        p_wishbone_bd_ram_n25023, p_wishbone_bd_ram_n25024, 
        p_wishbone_bd_ram_n25025, p_wishbone_bd_ram_n25026, 
        p_wishbone_bd_ram_n25027, p_wishbone_bd_ram_n25028, 
        p_wishbone_bd_ram_n25029, p_wishbone_bd_ram_n25030, 
        p_wishbone_bd_ram_n25031, p_wishbone_bd_ram_n25032, 
        p_wishbone_bd_ram_n25033, p_wishbone_bd_ram_n25034, 
        p_wishbone_bd_ram_n25035, p_wishbone_bd_ram_n25036, 
        p_wishbone_bd_ram_n25037, p_wishbone_bd_ram_n25038, 
        p_wishbone_bd_ram_n25039, p_wishbone_bd_ram_n25040, 
        p_wishbone_bd_ram_n25041, p_wishbone_bd_ram_n25042, 
        p_wishbone_bd_ram_n25043, p_wishbone_bd_ram_n25044, 
        p_wishbone_bd_ram_n25045, p_wishbone_bd_ram_n25046, 
        p_wishbone_bd_ram_n25047, p_wishbone_bd_ram_n25048, 
        p_wishbone_bd_ram_n25049, p_wishbone_bd_ram_n25050, 
        p_wishbone_bd_ram_n25051, p_wishbone_bd_ram_n25052, 
        p_wishbone_bd_ram_n25053, p_wishbone_bd_ram_n25054, 
        p_wishbone_bd_ram_n25055, p_wishbone_bd_ram_n25056, 
        p_wishbone_bd_ram_n25057, p_wishbone_bd_ram_n25058, 
        p_wishbone_bd_ram_n25059, p_wishbone_bd_ram_n25060, 
        p_wishbone_bd_ram_n25061, p_wishbone_bd_ram_n25062, 
        p_wishbone_bd_ram_n25063, p_wishbone_bd_ram_n25064, 
        p_wishbone_bd_ram_n25065, p_wishbone_bd_ram_n25066, 
        p_wishbone_bd_ram_n25067, p_wishbone_bd_ram_n25068, 
        p_wishbone_bd_ram_n25069, p_wishbone_bd_ram_n25070, 
        p_wishbone_bd_ram_n25071, p_wishbone_bd_ram_n25072, 
        p_wishbone_bd_ram_n25073, p_wishbone_bd_ram_n25074, 
        p_wishbone_bd_ram_n25075, p_wishbone_bd_ram_n25076, 
        p_wishbone_bd_ram_n25077, p_wishbone_bd_ram_n25078, 
        p_wishbone_bd_ram_n25079, p_wishbone_bd_ram_n25080, 
        p_wishbone_bd_ram_n25081, p_wishbone_bd_ram_n25082, 
        p_wishbone_bd_ram_n25083, p_wishbone_bd_ram_n25084, 
        p_wishbone_bd_ram_n25085, p_wishbone_bd_ram_n25086, 
        p_wishbone_bd_ram_n25087, p_wishbone_bd_ram_n25088, 
        p_wishbone_bd_ram_n25089, p_wishbone_bd_ram_n25090, 
        p_wishbone_bd_ram_n25091, p_wishbone_bd_ram_n25092, 
        p_wishbone_bd_ram_n25093, p_wishbone_bd_ram_n25094, 
        p_wishbone_bd_ram_n25095, p_wishbone_bd_ram_n25096, 
        p_wishbone_bd_ram_n25097, p_wishbone_bd_ram_n25098, 
        p_wishbone_bd_ram_n25099, p_wishbone_bd_ram_n25100, 
        p_wishbone_bd_ram_n25101, p_wishbone_bd_ram_n25102, 
        p_wishbone_bd_ram_n25103, p_wishbone_bd_ram_n25104, 
        p_wishbone_bd_ram_n25105, p_wishbone_bd_ram_n25106, 
        p_wishbone_bd_ram_n25107, p_wishbone_bd_ram_n25108, 
        p_wishbone_bd_ram_n25109, p_wishbone_bd_ram_n25110, 
        p_wishbone_bd_ram_n25111, p_wishbone_bd_ram_n25112, 
        p_wishbone_bd_ram_n25113, p_wishbone_bd_ram_n25114, 
        p_wishbone_bd_ram_n25115, p_wishbone_bd_ram_n25116, 
        p_wishbone_bd_ram_n25117, p_wishbone_bd_ram_n25118, 
        p_wishbone_bd_ram_n25119, p_wishbone_bd_ram_n25120, 
        p_wishbone_bd_ram_n25121, p_wishbone_bd_ram_n25122, 
        p_wishbone_bd_ram_n25123, p_wishbone_bd_ram_n25124, 
        p_wishbone_bd_ram_n25125, p_wishbone_bd_ram_n25126, 
        p_wishbone_bd_ram_n25127, p_wishbone_bd_ram_n25128, 
        p_wishbone_bd_ram_n25129, p_wishbone_bd_ram_n25130, 
        p_wishbone_bd_ram_n25131, p_wishbone_bd_ram_n25132, 
        p_wishbone_bd_ram_n25133, p_wishbone_bd_ram_n25134, 
        p_wishbone_bd_ram_n25135, p_wishbone_bd_ram_n25136, 
        p_wishbone_bd_ram_n25137, p_wishbone_bd_ram_n25138, 
        p_wishbone_bd_ram_n25139, p_wishbone_bd_ram_n25140, 
        p_wishbone_bd_ram_n25141, p_wishbone_bd_ram_n25142, 
        p_wishbone_bd_ram_n25143, p_wishbone_bd_ram_n25144, 
        p_wishbone_bd_ram_n25145, p_wishbone_bd_ram_n25146, 
        p_wishbone_bd_ram_n25147, p_wishbone_bd_ram_n25148, 
        p_wishbone_bd_ram_n25149, p_wishbone_bd_ram_n25150, 
        p_wishbone_bd_ram_n25151, p_wishbone_bd_ram_n25152, 
        p_wishbone_bd_ram_n25153, p_wishbone_bd_ram_n25154, 
        p_wishbone_bd_ram_n25155, p_wishbone_bd_ram_n25156, 
        p_wishbone_bd_ram_n25157, p_wishbone_bd_ram_n25158, 
        p_wishbone_bd_ram_n25159, p_wishbone_bd_ram_n25160, 
        p_wishbone_bd_ram_n25161, p_wishbone_bd_ram_n25162, 
        p_wishbone_bd_ram_n25163, p_wishbone_bd_ram_n25164, 
        p_wishbone_bd_ram_n25165, p_wishbone_bd_ram_n25166, 
        p_wishbone_bd_ram_n25167, p_wishbone_bd_ram_n25168, 
        p_wishbone_bd_ram_n25169, p_wishbone_bd_ram_n25170, 
        p_wishbone_bd_ram_n25171, p_wishbone_bd_ram_n25172, 
        p_wishbone_bd_ram_n25173, p_wishbone_bd_ram_n25174, 
        p_wishbone_bd_ram_n25175, p_wishbone_bd_ram_n25176, 
        p_wishbone_bd_ram_n25177, p_wishbone_bd_ram_n25178, 
        p_wishbone_bd_ram_n25179, p_wishbone_bd_ram_n25180, 
        p_wishbone_bd_ram_n25181, p_wishbone_bd_ram_n25182, 
        p_wishbone_bd_ram_n25183, p_wishbone_bd_ram_n25184, 
        p_wishbone_bd_ram_n25185, p_wishbone_bd_ram_n25186, 
        p_wishbone_bd_ram_n25187, p_wishbone_bd_ram_n25188, 
        p_wishbone_bd_ram_n25189, p_wishbone_bd_ram_n25190, 
        p_wishbone_bd_ram_n25191, p_wishbone_bd_ram_n25192, 
        p_wishbone_bd_ram_n25193, p_wishbone_bd_ram_n25194, 
        p_wishbone_bd_ram_n25195, p_wishbone_bd_ram_n25196, 
        p_wishbone_bd_ram_n25197, p_wishbone_bd_ram_n25198, 
        p_wishbone_bd_ram_n25199, p_wishbone_bd_ram_n25200, 
        p_wishbone_bd_ram_n25201, p_wishbone_bd_ram_n25202, 
        p_wishbone_bd_ram_n25203, p_wishbone_bd_ram_n25204, 
        p_wishbone_bd_ram_n25205, p_wishbone_bd_ram_n25206, 
        p_wishbone_bd_ram_n25207, p_wishbone_bd_ram_n25208, 
        p_wishbone_bd_ram_n25209, p_wishbone_bd_ram_n25210, 
        p_wishbone_bd_ram_n25211, p_wishbone_bd_ram_n25212, 
        p_wishbone_bd_ram_n25213, p_wishbone_bd_ram_n25214, 
        p_wishbone_bd_ram_n25215, p_wishbone_bd_ram_n25216, 
        p_wishbone_bd_ram_n25217, p_wishbone_bd_ram_n25218, 
        p_wishbone_bd_ram_n25219, p_wishbone_bd_ram_n25220, 
        p_wishbone_bd_ram_n25221, p_wishbone_bd_ram_n25222, 
        p_wishbone_bd_ram_n25223, p_wishbone_bd_ram_n25224, 
        p_wishbone_bd_ram_n25225, p_wishbone_bd_ram_n25226, 
        p_wishbone_bd_ram_n25227, p_wishbone_bd_ram_n25228, 
        p_wishbone_bd_ram_n25229, p_wishbone_bd_ram_n25230, 
        p_wishbone_bd_ram_n25231, p_wishbone_bd_ram_n25232, 
        p_wishbone_bd_ram_n25233, p_wishbone_bd_ram_n25234, 
        p_wishbone_bd_ram_n25235, p_wishbone_bd_ram_n25236, 
        p_wishbone_bd_ram_n25237, p_wishbone_bd_ram_n25238, 
        p_wishbone_bd_ram_n25239, p_wishbone_bd_ram_n25240, 
        p_wishbone_bd_ram_n25241, p_wishbone_bd_ram_n25242, 
        p_wishbone_bd_ram_n25243, p_wishbone_bd_ram_n25244, 
        p_wishbone_bd_ram_n25245, p_wishbone_bd_ram_n25246, 
        p_wishbone_bd_ram_n25247, p_wishbone_bd_ram_n25248, 
        p_wishbone_bd_ram_n25249, p_wishbone_bd_ram_n25250, 
        p_wishbone_bd_ram_n25251, p_wishbone_bd_ram_n25252, 
        p_wishbone_bd_ram_n25253, p_wishbone_bd_ram_n25254, 
        p_wishbone_bd_ram_n25255, p_wishbone_bd_ram_n25256, 
        p_wishbone_bd_ram_n25257, p_wishbone_bd_ram_n25258, 
        p_wishbone_bd_ram_n25259, p_wishbone_bd_ram_n25260, 
        p_wishbone_bd_ram_n25261, p_wishbone_bd_ram_n25262, 
        p_wishbone_bd_ram_n25263, p_wishbone_bd_ram_n25264, 
        p_wishbone_bd_ram_n25265, p_wishbone_bd_ram_n25266, 
        p_wishbone_bd_ram_n25267, p_wishbone_bd_ram_n25268, 
        p_wishbone_bd_ram_n25269, p_wishbone_bd_ram_n25270, 
        p_wishbone_bd_ram_n25271, p_wishbone_bd_ram_n25272, 
        p_wishbone_bd_ram_n25273, p_wishbone_bd_ram_n25274, 
        p_wishbone_bd_ram_n25275, p_wishbone_bd_ram_n25276, 
        p_wishbone_bd_ram_n25277, p_wishbone_bd_ram_n25278, 
        p_wishbone_bd_ram_n25279, p_wishbone_bd_ram_n25280, 
        p_wishbone_bd_ram_n25281, p_wishbone_bd_ram_n25282, 
        p_wishbone_bd_ram_n25283, p_wishbone_bd_ram_n25284, 
        p_wishbone_bd_ram_n25285, p_wishbone_bd_ram_n25286, 
        p_wishbone_bd_ram_n25287, p_wishbone_bd_ram_n25288, 
        p_wishbone_bd_ram_n25289, p_wishbone_bd_ram_n25290, 
        p_wishbone_bd_ram_n25291, p_wishbone_bd_ram_n25292, 
        p_wishbone_bd_ram_n25293, p_wishbone_bd_ram_n25294, 
        p_wishbone_bd_ram_n25295, p_wishbone_bd_ram_n25296, 
        p_wishbone_bd_ram_n25297, p_wishbone_bd_ram_n25298, 
        p_wishbone_bd_ram_n25299, p_wishbone_bd_ram_n25300, 
        p_wishbone_bd_ram_n25301, p_wishbone_bd_ram_n25302, 
        p_wishbone_bd_ram_n25303, p_wishbone_bd_ram_n25304, 
        p_wishbone_bd_ram_n25305, p_wishbone_bd_ram_n25306, 
        p_wishbone_bd_ram_n25307, p_wishbone_bd_ram_n25308, 
        p_wishbone_bd_ram_n25309, p_wishbone_bd_ram_n25310, 
        p_wishbone_bd_ram_n25311, p_wishbone_bd_ram_n25312, 
        p_wishbone_bd_ram_n25313, p_wishbone_bd_ram_n25314, 
        p_wishbone_bd_ram_n25315, p_wishbone_bd_ram_n25316, 
        p_wishbone_bd_ram_n25317, p_wishbone_bd_ram_n25318, 
        p_wishbone_bd_ram_n25319, p_wishbone_bd_ram_n25320, 
        p_wishbone_bd_ram_n25321, p_wishbone_bd_ram_n25322, 
        p_wishbone_bd_ram_n25323, p_wishbone_bd_ram_n25324, 
        p_wishbone_bd_ram_n25325, p_wishbone_bd_ram_n25326, 
        p_wishbone_bd_ram_n25327, p_wishbone_bd_ram_n25328, 
        p_wishbone_bd_ram_n25329, p_wishbone_bd_ram_n25330, 
        p_wishbone_bd_ram_n25331, p_wishbone_bd_ram_n25332, 
        p_wishbone_bd_ram_n25333, p_wishbone_bd_ram_n25334, 
        p_wishbone_bd_ram_n25335, p_wishbone_bd_ram_n25336, 
        p_wishbone_bd_ram_n25337, p_wishbone_bd_ram_n25338, 
        p_wishbone_bd_ram_n25339, p_wishbone_bd_ram_n25340, 
        p_wishbone_bd_ram_n25341, p_wishbone_bd_ram_n25342, 
        p_wishbone_bd_ram_n25343, p_wishbone_bd_ram_n25344, 
        p_wishbone_bd_ram_n25345, p_wishbone_bd_ram_n25346, 
        p_wishbone_bd_ram_n25347, p_wishbone_bd_ram_n25348, 
        p_wishbone_bd_ram_n25349, p_wishbone_bd_ram_n25350, 
        p_wishbone_bd_ram_n25351, p_wishbone_bd_ram_n25352, 
        p_wishbone_bd_ram_n25353, p_wishbone_bd_ram_n25354, 
        p_wishbone_bd_ram_n25355, p_wishbone_bd_ram_n25356, 
        p_wishbone_bd_ram_n25357, p_wishbone_bd_ram_n25358, 
        p_wishbone_bd_ram_n25359, p_wishbone_bd_ram_n25360, 
        p_wishbone_bd_ram_n25361, p_wishbone_bd_ram_n25362, 
        p_wishbone_bd_ram_n25363, p_wishbone_bd_ram_n25364, 
        p_wishbone_bd_ram_n25365, p_wishbone_bd_ram_n25366, 
        p_wishbone_bd_ram_n25367, p_wishbone_bd_ram_n25368, 
        p_wishbone_bd_ram_n25369, p_wishbone_bd_ram_n25370, 
        p_wishbone_bd_ram_n25371, p_wishbone_bd_ram_n25372, 
        p_wishbone_bd_ram_n25373, p_wishbone_bd_ram_n25374, 
        p_wishbone_bd_ram_n25375, p_wishbone_bd_ram_n25376, 
        p_wishbone_bd_ram_n25377, p_wishbone_bd_ram_n25378, 
        p_wishbone_bd_ram_n25379, p_wishbone_bd_ram_n25380, 
        p_wishbone_bd_ram_n25381, p_wishbone_bd_ram_n25382, 
        p_wishbone_bd_ram_n25383, p_wishbone_bd_ram_n25384, 
        p_wishbone_bd_ram_n25385, p_wishbone_bd_ram_n25386, 
        p_wishbone_bd_ram_n25387, p_wishbone_bd_ram_n25388, 
        p_wishbone_bd_ram_n25389, p_wishbone_bd_ram_n25390, 
        p_wishbone_bd_ram_n25391, p_wishbone_bd_ram_n25392, 
        p_wishbone_bd_ram_n25393, p_wishbone_bd_ram_n25394, 
        p_wishbone_bd_ram_n25395, p_wishbone_bd_ram_n25396, 
        p_wishbone_bd_ram_n25397, p_wishbone_bd_ram_n25398, 
        p_wishbone_bd_ram_n25399, p_wishbone_bd_ram_n25400, 
        p_wishbone_bd_ram_n25401, p_wishbone_bd_ram_n25402, 
        p_wishbone_bd_ram_n25403, p_wishbone_bd_ram_n25404, 
        p_wishbone_bd_ram_n25405, p_wishbone_bd_ram_n25406, 
        p_wishbone_bd_ram_n25407, p_wishbone_bd_ram_n25408, 
        p_wishbone_bd_ram_n25409, p_wishbone_bd_ram_n25410, 
        p_wishbone_bd_ram_n25411, p_wishbone_bd_ram_n25412, 
        p_wishbone_bd_ram_n25413, p_wishbone_bd_ram_n25414, 
        p_wishbone_bd_ram_n25415, p_wishbone_bd_ram_n25416, 
        p_wishbone_bd_ram_n25417, p_wishbone_bd_ram_n25418, 
        p_wishbone_bd_ram_n25419, p_wishbone_bd_ram_n25420, 
        p_wishbone_bd_ram_n25421, p_wishbone_bd_ram_n25422, 
        p_wishbone_bd_ram_n25423, p_wishbone_bd_ram_n25424, 
        p_wishbone_bd_ram_n25425, p_wishbone_bd_ram_n25426, 
        p_wishbone_bd_ram_n25427, p_wishbone_bd_ram_n25428, 
        p_wishbone_bd_ram_n25429, p_wishbone_bd_ram_n25430, 
        p_wishbone_bd_ram_n25431, p_wishbone_bd_ram_n25432, 
        p_wishbone_bd_ram_n25433, p_wishbone_bd_ram_n25434, 
        p_wishbone_bd_ram_n25435, p_wishbone_bd_ram_n25436, 
        p_wishbone_bd_ram_n25437, p_wishbone_bd_ram_n25438, 
        p_wishbone_bd_ram_n25439, p_wishbone_bd_ram_n25440, 
        p_wishbone_bd_ram_n25441, p_wishbone_bd_ram_n25442, 
        p_wishbone_bd_ram_n25443, p_wishbone_bd_ram_n25444, 
        p_wishbone_bd_ram_n25445, p_wishbone_bd_ram_n25446, 
        p_wishbone_bd_ram_n25447, p_wishbone_bd_ram_n25448, 
        p_wishbone_bd_ram_n25449, p_wishbone_bd_ram_n25450, 
        p_wishbone_bd_ram_n25451, p_wishbone_bd_ram_n25452, 
        p_wishbone_bd_ram_n25453, p_wishbone_bd_ram_n25454, 
        p_wishbone_bd_ram_n25455, p_wishbone_bd_ram_n25456, 
        p_wishbone_bd_ram_n25457, p_wishbone_bd_ram_n25458, 
        p_wishbone_bd_ram_n25459, p_wishbone_bd_ram_n25460, 
        p_wishbone_bd_ram_n25461, p_wishbone_bd_ram_n25462, 
        p_wishbone_bd_ram_n25463, p_wishbone_bd_ram_n25464, 
        p_wishbone_bd_ram_n25465, p_wishbone_bd_ram_n25466, 
        p_wishbone_bd_ram_n25467, p_wishbone_bd_ram_n25468, 
        p_wishbone_bd_ram_n25469, p_wishbone_bd_ram_n25470, 
        p_wishbone_bd_ram_n25471, p_wishbone_bd_ram_n25472, 
        p_wishbone_bd_ram_n25473, p_wishbone_bd_ram_n25474, 
        p_wishbone_bd_ram_n25475, p_wishbone_bd_ram_n25476, 
        p_wishbone_bd_ram_n25477, p_wishbone_bd_ram_n25478, 
        p_wishbone_bd_ram_n25479, p_wishbone_bd_ram_n25480, 
        p_wishbone_bd_ram_n25481, p_wishbone_bd_ram_n25482, 
        p_wishbone_bd_ram_n25483, p_wishbone_bd_ram_n25484, 
        p_wishbone_bd_ram_n25485, p_wishbone_bd_ram_n25486, 
        p_wishbone_bd_ram_n25487, p_wishbone_bd_ram_n25488, 
        p_wishbone_bd_ram_n25489, p_wishbone_bd_ram_n25490, 
        p_wishbone_bd_ram_n25491, p_wishbone_bd_ram_n25492, 
        p_wishbone_bd_ram_n25493, p_wishbone_bd_ram_n25494, 
        p_wishbone_bd_ram_n25495, p_wishbone_bd_ram_n25496, 
        p_wishbone_bd_ram_n25497, p_wishbone_bd_ram_n25498, 
        p_wishbone_bd_ram_n25499, p_wishbone_bd_ram_n25500, 
        p_wishbone_bd_ram_n25501, p_wishbone_bd_ram_n25502, 
        p_wishbone_bd_ram_n25503, p_wishbone_bd_ram_n25504, 
        p_wishbone_bd_ram_n25505, p_wishbone_bd_ram_n25506, 
        p_wishbone_bd_ram_n25507, p_wishbone_bd_ram_n25508, 
        p_wishbone_bd_ram_n25509, p_wishbone_bd_ram_n25510, 
        p_wishbone_bd_ram_n25511, p_wishbone_bd_ram_n25512, 
        p_wishbone_bd_ram_n25513, p_wishbone_bd_ram_n25514, 
        p_wishbone_bd_ram_n25515, p_wishbone_bd_ram_n25516, 
        p_wishbone_bd_ram_n25517, p_wishbone_bd_ram_n25518, 
        p_wishbone_bd_ram_n25519, p_wishbone_bd_ram_n25520, 
        p_wishbone_bd_ram_n25521, p_wishbone_bd_ram_n25522, 
        p_wishbone_bd_ram_n25523, p_wishbone_bd_ram_n25524, 
        p_wishbone_bd_ram_n25525, p_wishbone_bd_ram_n25526, 
        p_wishbone_bd_ram_n25527, p_wishbone_bd_ram_n25528, 
        p_wishbone_bd_ram_n25529, p_wishbone_bd_ram_n25530, 
        p_wishbone_bd_ram_n25531, p_wishbone_bd_ram_n25532, 
        p_wishbone_bd_ram_n25533, p_wishbone_bd_ram_n25534, 
        p_wishbone_bd_ram_n25535, p_wishbone_bd_ram_n25536, 
        p_wishbone_bd_ram_n25537, p_wishbone_bd_ram_n25538, 
        p_wishbone_bd_ram_n25539, p_wishbone_bd_ram_n25540, 
        p_wishbone_bd_ram_n25541, p_wishbone_bd_ram_n25542, 
        p_wishbone_bd_ram_n25543, p_wishbone_bd_ram_n25544, 
        p_wishbone_bd_ram_n25545, p_wishbone_bd_ram_n25546, 
        p_wishbone_bd_ram_n25547, p_wishbone_bd_ram_n25548, 
        p_wishbone_bd_ram_n25549, p_wishbone_bd_ram_n25550, 
        p_wishbone_bd_ram_n25551, p_wishbone_bd_ram_n25552, 
        p_wishbone_bd_ram_n25553, p_wishbone_bd_ram_n25554, 
        p_wishbone_bd_ram_n25555, p_wishbone_bd_ram_n25556, 
        p_wishbone_bd_ram_n25557, p_wishbone_bd_ram_n25558, 
        p_wishbone_bd_ram_n25559, p_wishbone_bd_ram_n25560, 
        p_wishbone_bd_ram_n25561, p_wishbone_bd_ram_n25562, 
        p_wishbone_bd_ram_n25563, p_wishbone_bd_ram_n25564, 
        p_wishbone_bd_ram_n25565, p_wishbone_bd_ram_n25566, 
        p_wishbone_bd_ram_n25567, p_wishbone_bd_ram_n25568, 
        p_wishbone_bd_ram_n25569, p_wishbone_bd_ram_n25570, 
        p_wishbone_bd_ram_n25571, p_wishbone_bd_ram_n25572, 
        p_wishbone_bd_ram_n25573, p_wishbone_bd_ram_n25574, 
        p_wishbone_bd_ram_n25575, p_wishbone_bd_ram_n25576, 
        p_wishbone_bd_ram_n25577, p_wishbone_bd_ram_n25578, 
        p_wishbone_bd_ram_n25579, p_wishbone_bd_ram_n25580, 
        p_wishbone_bd_ram_n25581, p_wishbone_bd_ram_n25582, 
        p_wishbone_bd_ram_n25583, p_wishbone_bd_ram_n25584, 
        p_wishbone_bd_ram_n25585, p_wishbone_bd_ram_n25586, 
        p_wishbone_bd_ram_n25587, p_wishbone_bd_ram_n25588, 
        p_wishbone_bd_ram_n25589, p_wishbone_bd_ram_n25590, 
        p_wishbone_bd_ram_n25591, p_wishbone_bd_ram_n25592, 
        p_wishbone_bd_ram_n25593, p_wishbone_bd_ram_n25594, 
        p_wishbone_bd_ram_n25595, p_wishbone_bd_ram_n25596, 
        p_wishbone_bd_ram_n25597, p_wishbone_bd_ram_n25598, 
        p_wishbone_bd_ram_n25599, p_wishbone_bd_ram_n25600, 
        p_wishbone_bd_ram_n25601, p_wishbone_bd_ram_n25602, 
        p_wishbone_bd_ram_n25603, p_wishbone_bd_ram_n25604, 
        p_wishbone_bd_ram_n25605, p_wishbone_bd_ram_n25606, 
        p_wishbone_bd_ram_n25607, p_wishbone_bd_ram_n25608, 
        p_wishbone_bd_ram_n25609, p_wishbone_bd_ram_n25610, 
        p_wishbone_bd_ram_n25611, p_wishbone_bd_ram_n25612, 
        p_wishbone_bd_ram_n25613, p_wishbone_bd_ram_n25614, 
        p_wishbone_bd_ram_n25615, p_wishbone_bd_ram_n25616, 
        p_wishbone_bd_ram_n25617, p_wishbone_bd_ram_n25618, 
        p_wishbone_bd_ram_n25619, p_wishbone_bd_ram_n25620, 
        p_wishbone_bd_ram_n25621, p_wishbone_bd_ram_n25622, 
        p_wishbone_bd_ram_n25623, p_wishbone_bd_ram_n25624, 
        p_wishbone_bd_ram_n25625, p_wishbone_bd_ram_n25626, 
        p_wishbone_bd_ram_n25627, p_wishbone_bd_ram_n25628, 
        p_wishbone_bd_ram_n25629, p_wishbone_bd_ram_n25630, 
        p_wishbone_bd_ram_n25631, p_wishbone_bd_ram_n25632, 
        p_wishbone_bd_ram_n25633, p_wishbone_bd_ram_n25634, 
        p_wishbone_bd_ram_n25635, p_wishbone_bd_ram_n25636, 
        p_wishbone_bd_ram_n25637, p_wishbone_bd_ram_n25638, 
        p_wishbone_bd_ram_n25639, p_wishbone_bd_ram_n25640, 
        p_wishbone_bd_ram_n25641, p_wishbone_bd_ram_n25642, 
        p_wishbone_bd_ram_n25643, p_wishbone_bd_ram_n25644, 
        p_wishbone_bd_ram_n25645, p_wishbone_bd_ram_n25646, 
        p_wishbone_bd_ram_n25647, p_wishbone_bd_ram_n25648, 
        p_wishbone_bd_ram_n25649, p_wishbone_bd_ram_n25650, 
        p_wishbone_bd_ram_n25651, p_wishbone_bd_ram_n25652, 
        p_wishbone_bd_ram_n25653, p_wishbone_bd_ram_n25654, 
        p_wishbone_bd_ram_n25655, p_wishbone_bd_ram_n25656, 
        p_wishbone_bd_ram_n25657, p_wishbone_bd_ram_n25658, 
        p_wishbone_bd_ram_n25659, p_wishbone_bd_ram_n25660, 
        p_wishbone_bd_ram_n25661, p_wishbone_bd_ram_n25662, 
        p_wishbone_bd_ram_n25663, p_wishbone_bd_ram_n25664, 
        p_wishbone_bd_ram_n25665, p_wishbone_bd_ram_n25666, 
        p_wishbone_bd_ram_n25667, p_wishbone_bd_ram_n25668, 
        p_wishbone_bd_ram_n25669, p_wishbone_bd_ram_n25670, 
        p_wishbone_bd_ram_n25671, p_wishbone_bd_ram_n25672, 
        p_wishbone_bd_ram_n25673, p_wishbone_bd_ram_n25674, 
        p_wishbone_bd_ram_n25675, p_wishbone_bd_ram_n25676, 
        p_wishbone_bd_ram_n25677, p_wishbone_bd_ram_n25678, 
        p_wishbone_bd_ram_n25679, p_wishbone_bd_ram_n25680, 
        p_wishbone_bd_ram_n25681, p_wishbone_bd_ram_n25682, 
        p_wishbone_bd_ram_n25683, p_wishbone_bd_ram_n25684, 
        p_wishbone_bd_ram_n25685, p_wishbone_bd_ram_n25686, 
        p_wishbone_bd_ram_n25687, p_wishbone_bd_ram_n25688, 
        p_wishbone_bd_ram_n25689, p_wishbone_bd_ram_n25690, 
        p_wishbone_bd_ram_n25691, p_wishbone_bd_ram_n25692, 
        p_wishbone_bd_ram_n25693, p_wishbone_bd_ram_n25694, 
        p_wishbone_bd_ram_n25695, p_wishbone_bd_ram_n25696, 
        p_wishbone_bd_ram_n25697, p_wishbone_bd_ram_n25698, 
        p_wishbone_bd_ram_n25699, p_wishbone_bd_ram_n25700, 
        p_wishbone_bd_ram_n25701, p_wishbone_bd_ram_n25702, 
        p_wishbone_bd_ram_n25703, p_wishbone_bd_ram_n25704, 
        p_wishbone_bd_ram_n25705, p_wishbone_bd_ram_n25706, 
        p_wishbone_bd_ram_n25707, p_wishbone_bd_ram_n25708, 
        p_wishbone_bd_ram_n25709, p_wishbone_bd_ram_n25710, 
        p_wishbone_bd_ram_n25711, p_wishbone_bd_ram_n25712, 
        p_wishbone_bd_ram_n25713, p_wishbone_bd_ram_n25714, 
        p_wishbone_bd_ram_n25715, p_wishbone_bd_ram_n25716, 
        p_wishbone_bd_ram_n25717, p_wishbone_bd_ram_n25718, 
        p_wishbone_bd_ram_n25719, p_wishbone_bd_ram_n25720, 
        p_wishbone_bd_ram_n25721, p_wishbone_bd_ram_n25722, 
        p_wishbone_bd_ram_n25723, p_wishbone_bd_ram_n25724, 
        p_wishbone_bd_ram_n25725, p_wishbone_bd_ram_n25726, 
        p_wishbone_bd_ram_n25727, p_wishbone_bd_ram_n25728, 
        p_wishbone_bd_ram_n25729, p_wishbone_bd_ram_n25730, 
        p_wishbone_bd_ram_n25731, p_wishbone_bd_ram_n25732, 
        p_wishbone_bd_ram_n25733, p_wishbone_bd_ram_n25734, 
        p_wishbone_bd_ram_n25735, p_wishbone_bd_ram_n25736, 
        p_wishbone_bd_ram_n25737, p_wishbone_bd_ram_n25738, 
        p_wishbone_bd_ram_n25739, p_wishbone_bd_ram_n25740, 
        p_wishbone_bd_ram_n25741, p_wishbone_bd_ram_n25742, 
        p_wishbone_bd_ram_n25743, p_wishbone_bd_ram_n25744, 
        p_wishbone_bd_ram_n25745, p_wishbone_bd_ram_n25746, 
        p_wishbone_bd_ram_n25747, p_wishbone_bd_ram_n25748, 
        p_wishbone_bd_ram_n25749, p_wishbone_bd_ram_n25750, 
        p_wishbone_bd_ram_n25751, p_wishbone_bd_ram_n25752, 
        p_wishbone_bd_ram_n25753, p_wishbone_bd_ram_n25754, 
        p_wishbone_bd_ram_n25755, p_wishbone_bd_ram_n25756, 
        p_wishbone_bd_ram_n25757, p_wishbone_bd_ram_n25758, 
        p_wishbone_bd_ram_n25759, p_wishbone_bd_ram_n25760, 
        p_wishbone_bd_ram_n25761, p_wishbone_bd_ram_n25762, 
        p_wishbone_bd_ram_n25763, p_wishbone_bd_ram_n25764, 
        p_wishbone_bd_ram_n25765, p_wishbone_bd_ram_n25766, 
        p_wishbone_bd_ram_n25767, p_wishbone_bd_ram_n25768, 
        p_wishbone_bd_ram_n25769, p_wishbone_bd_ram_n25770, 
        p_wishbone_bd_ram_n25771, p_wishbone_bd_ram_n25772, 
        p_wishbone_bd_ram_n25773, p_wishbone_bd_ram_n25774, 
        p_wishbone_bd_ram_n25775, p_wishbone_bd_ram_n25776, 
        p_wishbone_bd_ram_n25777, p_wishbone_bd_ram_n25778, 
        p_wishbone_bd_ram_n25779, p_wishbone_bd_ram_n25780, 
        p_wishbone_bd_ram_n25781, p_wishbone_bd_ram_n25782, 
        p_wishbone_bd_ram_n25783, p_wishbone_bd_ram_n25784, 
        p_wishbone_bd_ram_n25785, p_wishbone_bd_ram_n25786, 
        p_wishbone_bd_ram_n25787, p_wishbone_bd_ram_n25788, 
        p_wishbone_bd_ram_n25789, p_wishbone_bd_ram_n25790, 
        p_wishbone_bd_ram_n25791, p_wishbone_bd_ram_n25792, 
        p_wishbone_bd_ram_n25793, p_wishbone_bd_ram_n25794, 
        p_wishbone_bd_ram_n25795, p_wishbone_bd_ram_n25796, 
        p_wishbone_bd_ram_n25797, p_wishbone_bd_ram_n25798, 
        p_wishbone_bd_ram_n25799, p_wishbone_bd_ram_n25800, 
        p_wishbone_bd_ram_n25801, p_wishbone_bd_ram_n25802, 
        p_wishbone_bd_ram_n25803, p_wishbone_bd_ram_n25804, 
        p_wishbone_bd_ram_n25805, p_wishbone_bd_ram_n25806, 
        p_wishbone_bd_ram_n25807, p_wishbone_bd_ram_n25808, 
        p_wishbone_bd_ram_n25809, p_wishbone_bd_ram_n25810, 
        p_wishbone_bd_ram_n25811, p_wishbone_bd_ram_n25812, 
        p_wishbone_bd_ram_n25813, p_wishbone_bd_ram_n25814, 
        p_wishbone_bd_ram_n25815, p_wishbone_bd_ram_n25816, 
        p_wishbone_bd_ram_n25817, p_wishbone_bd_ram_n25818, 
        p_wishbone_bd_ram_n25819, p_wishbone_bd_ram_n25820, 
        p_wishbone_bd_ram_n25821, p_wishbone_bd_ram_n25822, 
        p_wishbone_bd_ram_n25823, p_wishbone_bd_ram_n25824, 
        p_wishbone_bd_ram_n25825, p_wishbone_bd_ram_n25826, 
        p_wishbone_bd_ram_n25827, p_wishbone_bd_ram_n25828, 
        p_wishbone_bd_ram_n25829, p_wishbone_bd_ram_n25830, 
        p_wishbone_bd_ram_n25831, p_wishbone_bd_ram_n25832, 
        p_wishbone_bd_ram_n25833, p_wishbone_bd_ram_n25834, 
        p_wishbone_bd_ram_n25835, p_wishbone_bd_ram_n25836, 
        p_wishbone_bd_ram_n25837, p_wishbone_bd_ram_n25838, 
        p_wishbone_bd_ram_n25839, p_wishbone_bd_ram_n25840, 
        p_wishbone_bd_ram_n25841, p_wishbone_bd_ram_n25842, 
        p_wishbone_bd_ram_n25843, p_wishbone_bd_ram_n25844, 
        p_wishbone_bd_ram_n25845, p_wishbone_bd_ram_n25846, 
        p_wishbone_bd_ram_n25847, p_wishbone_bd_ram_n25848, 
        p_wishbone_bd_ram_n25849, p_wishbone_bd_ram_n25850, 
        p_wishbone_bd_ram_n25851, p_wishbone_bd_ram_n25852, 
        p_wishbone_bd_ram_n25853, p_wishbone_bd_ram_n25854, 
        p_wishbone_bd_ram_n25855, p_wishbone_bd_ram_n25856, 
        p_wishbone_bd_ram_n25857, p_wishbone_bd_ram_n25858, 
        p_wishbone_bd_ram_n25859, p_wishbone_bd_ram_n25860, 
        p_wishbone_bd_ram_n25861, p_wishbone_bd_ram_n25862, 
        p_wishbone_bd_ram_n25863, p_wishbone_bd_ram_n25864, 
        p_wishbone_bd_ram_n25865, p_wishbone_bd_ram_n25866, 
        p_wishbone_bd_ram_n25867, p_wishbone_bd_ram_n25868, 
        p_wishbone_bd_ram_n25869, p_wishbone_bd_ram_n25870, 
        p_wishbone_bd_ram_n25871, p_wishbone_bd_ram_n25872, 
        p_wishbone_bd_ram_n25873, p_wishbone_bd_ram_n25874, 
        p_wishbone_bd_ram_n25875, p_wishbone_bd_ram_n25876, 
        p_wishbone_bd_ram_n25877, p_wishbone_bd_ram_n25878, 
        p_wishbone_bd_ram_n25879, p_wishbone_bd_ram_n25880, 
        p_wishbone_bd_ram_n25881, p_wishbone_bd_ram_n25882, 
        p_wishbone_bd_ram_n25883, p_wishbone_bd_ram_n25884, 
        p_wishbone_bd_ram_n25885, p_wishbone_bd_ram_n25886, 
        p_wishbone_bd_ram_n25887, p_wishbone_bd_ram_n25888, 
        p_wishbone_bd_ram_n25889, p_wishbone_bd_ram_n25890, 
        p_wishbone_bd_ram_n25891, p_wishbone_bd_ram_n25892, 
        p_wishbone_bd_ram_n25893, p_wishbone_bd_ram_n25894, 
        p_wishbone_bd_ram_n25895, p_wishbone_bd_ram_n25896, 
        p_wishbone_bd_ram_n25897, p_wishbone_bd_ram_n25898, 
        p_wishbone_bd_ram_n25899, p_wishbone_bd_ram_n25900, 
        p_wishbone_bd_ram_n25901, p_wishbone_bd_ram_n25902, 
        p_wishbone_bd_ram_n25903, p_wishbone_bd_ram_n25904, 
        p_wishbone_bd_ram_n25905, p_wishbone_bd_ram_n25906, 
        p_wishbone_bd_ram_n25907, p_wishbone_bd_ram_n25908, 
        p_wishbone_bd_ram_n25909, p_wishbone_bd_ram_n25910, 
        p_wishbone_bd_ram_n25911, p_wishbone_bd_ram_n25912, 
        p_wishbone_bd_ram_n25913, p_wishbone_bd_ram_n25914, 
        p_wishbone_bd_ram_n25915, p_wishbone_bd_ram_n25916, 
        p_wishbone_bd_ram_n25917, p_wishbone_bd_ram_n25918, 
        p_wishbone_bd_ram_n25919, p_wishbone_bd_ram_n25920, 
        p_wishbone_bd_ram_n25921, p_wishbone_bd_ram_n25922, 
        p_wishbone_bd_ram_n25923, p_wishbone_bd_ram_n25924, 
        p_wishbone_bd_ram_n25925, p_wishbone_bd_ram_n25926, 
        p_wishbone_bd_ram_n25927, p_wishbone_bd_ram_n25928, 
        p_wishbone_bd_ram_n25929, p_wishbone_bd_ram_n25930, 
        p_wishbone_bd_ram_n25931, p_wishbone_bd_ram_n25932, 
        p_wishbone_bd_ram_n25933, p_wishbone_bd_ram_n25934, 
        p_wishbone_bd_ram_n25935, p_wishbone_bd_ram_n25936, 
        p_wishbone_bd_ram_n25937, p_wishbone_bd_ram_n25938, 
        p_wishbone_bd_ram_n25939, p_wishbone_bd_ram_n25940, 
        p_wishbone_bd_ram_n25941, p_wishbone_bd_ram_n25942, 
        p_wishbone_bd_ram_n25943, p_wishbone_bd_ram_n25944, 
        p_wishbone_bd_ram_n25945, p_wishbone_bd_ram_n25946, 
        p_wishbone_bd_ram_n25947, p_wishbone_bd_ram_n25948, 
        p_wishbone_bd_ram_n25949, p_wishbone_bd_ram_n25950, 
        p_wishbone_bd_ram_n25951, p_wishbone_bd_ram_n25952, 
        p_wishbone_bd_ram_n25953, p_wishbone_bd_ram_n25954, 
        p_wishbone_bd_ram_n25955, p_wishbone_bd_ram_n25956, 
        p_wishbone_bd_ram_n25957, p_wishbone_bd_ram_n25958, 
        p_wishbone_bd_ram_n25959, p_wishbone_bd_ram_n25960, 
        p_wishbone_bd_ram_n25961, p_wishbone_bd_ram_n25962, 
        p_wishbone_bd_ram_n25963, p_wishbone_bd_ram_n25964, 
        p_wishbone_bd_ram_n25965, p_wishbone_bd_ram_n25966, 
        p_wishbone_bd_ram_n25967, p_wishbone_bd_ram_n25968, 
        p_wishbone_bd_ram_n25969, p_wishbone_bd_ram_n25970, 
        p_wishbone_bd_ram_n25971, p_wishbone_bd_ram_n25972, 
        p_wishbone_bd_ram_n25973, p_wishbone_bd_ram_n25974, 
        p_wishbone_bd_ram_n25975, p_wishbone_bd_ram_n25976, 
        p_wishbone_bd_ram_n25977, p_wishbone_bd_ram_n25978, 
        p_wishbone_bd_ram_n25979, p_wishbone_bd_ram_n25980, 
        p_wishbone_bd_ram_n25981, p_wishbone_bd_ram_n25982, 
        p_wishbone_bd_ram_n25983, p_wishbone_bd_ram_n25984, 
        p_wishbone_tx_fifo_N623, p_wishbone_tx_fifo_N624, 
        p_wishbone_tx_fifo_N625, p_wishbone_tx_fifo_N626, 
        p_wishbone_tx_fifo_N627, p_wishbone_tx_fifo_N628, 
        p_wishbone_tx_fifo_N629, p_wishbone_tx_fifo_N630, 
        p_wishbone_tx_fifo_N631, p_wishbone_tx_fifo_N632, 
        p_wishbone_tx_fifo_N633, p_wishbone_tx_fifo_N634, 
        p_wishbone_tx_fifo_N635, p_wishbone_tx_fifo_N636, 
        p_wishbone_tx_fifo_N637, p_wishbone_tx_fifo_N638, 
        p_wishbone_tx_fifo_N639, p_wishbone_tx_fifo_N640, 
        p_wishbone_tx_fifo_N641, p_wishbone_tx_fifo_N642, 
        p_wishbone_tx_fifo_N643, p_wishbone_tx_fifo_N644, 
        p_wishbone_tx_fifo_N645, p_wishbone_tx_fifo_N646, 
        p_wishbone_tx_fifo_N647, p_wishbone_tx_fifo_N648, 
        p_wishbone_tx_fifo_N649, p_wishbone_tx_fifo_N650, 
        p_wishbone_tx_fifo_N651, p_wishbone_tx_fifo_N652, 
        p_wishbone_tx_fifo_N653, p_wishbone_tx_fifo_N654, 
        p_wishbone_tx_fifo_n1229, p_wishbone_tx_fifo_n1230, 
        p_wishbone_tx_fifo_n1231, p_wishbone_tx_fifo_n1232, 
        p_wishbone_tx_fifo_n1233, p_wishbone_tx_fifo_n1234, 
        p_wishbone_tx_fifo_n1235, p_wishbone_tx_fifo_n1236, 
        p_wishbone_tx_fifo_n1237, p_wishbone_tx_fifo_n1238, 
        p_wishbone_tx_fifo_n1239, p_wishbone_tx_fifo_n1240, 
        p_wishbone_tx_fifo_n1241, p_wishbone_tx_fifo_n1242, 
        p_wishbone_tx_fifo_n1243, p_wishbone_tx_fifo_n1244, 
        p_wishbone_tx_fifo_n1245, p_wishbone_tx_fifo_n1246, 
        p_wishbone_tx_fifo_n1247, p_wishbone_tx_fifo_n1248, 
        p_wishbone_tx_fifo_n1249, p_wishbone_tx_fifo_n1250, 
        p_wishbone_tx_fifo_n1251, p_wishbone_tx_fifo_n1252, 
        p_wishbone_tx_fifo_n1253, p_wishbone_tx_fifo_n1254, 
        p_wishbone_tx_fifo_n1255, p_wishbone_tx_fifo_n1256, 
        p_wishbone_tx_fifo_n1257, p_wishbone_tx_fifo_n1258, 
        p_wishbone_tx_fifo_n1259, p_wishbone_tx_fifo_n1260, 
        p_wishbone_tx_fifo_n1261, p_wishbone_tx_fifo_n1262, 
        p_wishbone_tx_fifo_n1263, p_wishbone_tx_fifo_n1264, 
        p_wishbone_tx_fifo_n1265, p_wishbone_tx_fifo_n1266, 
        p_wishbone_tx_fifo_n1267, p_wishbone_tx_fifo_n1268, 
        p_wishbone_tx_fifo_n1269, p_wishbone_tx_fifo_n1270, 
        p_wishbone_tx_fifo_n1271, p_wishbone_tx_fifo_n1272, 
        p_wishbone_tx_fifo_n1273, p_wishbone_tx_fifo_n1274, 
        p_wishbone_tx_fifo_n1275, p_wishbone_tx_fifo_n1276, 
        p_wishbone_tx_fifo_n1277, p_wishbone_tx_fifo_n1278, 
        p_wishbone_tx_fifo_n1279, p_wishbone_tx_fifo_n1280, 
        p_wishbone_tx_fifo_n1281, p_wishbone_tx_fifo_n1282, 
        p_wishbone_tx_fifo_n1283, p_wishbone_tx_fifo_n1284, 
        p_wishbone_tx_fifo_n1285, p_wishbone_tx_fifo_n1286, 
        p_wishbone_tx_fifo_n1287, p_wishbone_tx_fifo_n1288, 
        p_wishbone_tx_fifo_n1289, p_wishbone_tx_fifo_n1290, 
        p_wishbone_tx_fifo_n1291, p_wishbone_tx_fifo_n1292, 
        p_wishbone_tx_fifo_n1293, p_wishbone_tx_fifo_n1294, 
        p_wishbone_tx_fifo_n1295, p_wishbone_tx_fifo_n1296, 
        p_wishbone_tx_fifo_n1297, p_wishbone_tx_fifo_n1298, 
        p_wishbone_tx_fifo_n1299, p_wishbone_tx_fifo_n1300, 
        p_wishbone_tx_fifo_n1301, p_wishbone_tx_fifo_n1302, 
        p_wishbone_tx_fifo_n1303, p_wishbone_tx_fifo_n1304, 
        p_wishbone_tx_fifo_n1305, p_wishbone_tx_fifo_n1306, 
        p_wishbone_tx_fifo_n1307, p_wishbone_tx_fifo_n1308, 
        p_wishbone_tx_fifo_n1309, p_wishbone_tx_fifo_n1310, 
        p_wishbone_tx_fifo_n1311, p_wishbone_tx_fifo_n1312, 
        p_wishbone_tx_fifo_n1313, p_wishbone_tx_fifo_n1314, 
        p_wishbone_tx_fifo_n1315, p_wishbone_tx_fifo_n1316, 
        p_wishbone_tx_fifo_n1317, p_wishbone_tx_fifo_n1318, 
        p_wishbone_tx_fifo_n1319, p_wishbone_tx_fifo_n1320, 
        p_wishbone_tx_fifo_n1321, p_wishbone_tx_fifo_n1322, 
        p_wishbone_tx_fifo_n1323, p_wishbone_tx_fifo_n1324, 
        p_wishbone_tx_fifo_n1325, p_wishbone_tx_fifo_n1326, 
        p_wishbone_tx_fifo_n1327, p_wishbone_tx_fifo_n1328, 
        p_wishbone_tx_fifo_n1329, p_wishbone_tx_fifo_n1330, 
        p_wishbone_tx_fifo_n1331, p_wishbone_tx_fifo_n1332, 
        p_wishbone_tx_fifo_n1333, p_wishbone_tx_fifo_n1334, 
        p_wishbone_tx_fifo_n1335, p_wishbone_tx_fifo_n1336, 
        p_wishbone_tx_fifo_n1337, p_wishbone_tx_fifo_n1338, 
        p_wishbone_tx_fifo_n1339, p_wishbone_tx_fifo_n1340, 
        p_wishbone_tx_fifo_n1341, p_wishbone_tx_fifo_n1342, 
        p_wishbone_tx_fifo_n1343, p_wishbone_tx_fifo_n1344, 
        p_wishbone_tx_fifo_n1345, p_wishbone_tx_fifo_n1346, 
        p_wishbone_tx_fifo_n1347, p_wishbone_tx_fifo_n1348, 
        p_wishbone_tx_fifo_n1349, p_wishbone_tx_fifo_n1350, 
        p_wishbone_tx_fifo_n1351, p_wishbone_tx_fifo_n1352, 
        p_wishbone_tx_fifo_n1353, p_wishbone_tx_fifo_n1354, 
        p_wishbone_tx_fifo_n1355, p_wishbone_tx_fifo_n1356, 
        p_wishbone_tx_fifo_n1357, p_wishbone_tx_fifo_n1358, 
        p_wishbone_tx_fifo_n1359, p_wishbone_tx_fifo_n1360, 
        p_wishbone_tx_fifo_n1361, p_wishbone_tx_fifo_n1362, 
        p_wishbone_tx_fifo_n1363, p_wishbone_tx_fifo_n1364, 
        p_wishbone_tx_fifo_n1365, p_wishbone_tx_fifo_n1366, 
        p_wishbone_tx_fifo_n1367, p_wishbone_tx_fifo_n1368, 
        p_wishbone_tx_fifo_n1369, p_wishbone_tx_fifo_n1370, 
        p_wishbone_tx_fifo_n1371, p_wishbone_tx_fifo_n1372, 
        p_wishbone_tx_fifo_n1373, p_wishbone_tx_fifo_n1374, 
        p_wishbone_tx_fifo_n1375, p_wishbone_tx_fifo_n1376, 
        p_wishbone_tx_fifo_n1377, p_wishbone_tx_fifo_n1378, 
        p_wishbone_tx_fifo_n1379, p_wishbone_tx_fifo_n1380, 
        p_wishbone_tx_fifo_n1381, p_wishbone_tx_fifo_n1382, 
        p_wishbone_tx_fifo_n1383, p_wishbone_tx_fifo_n1384, 
        p_wishbone_tx_fifo_n1385, p_wishbone_tx_fifo_n1386, 
        p_wishbone_tx_fifo_n1387, p_wishbone_tx_fifo_n1388, 
        p_wishbone_tx_fifo_n1389, p_wishbone_tx_fifo_n1390, 
        p_wishbone_tx_fifo_n1391, p_wishbone_tx_fifo_n1392, 
        p_wishbone_tx_fifo_n1393, p_wishbone_tx_fifo_n1394, 
        p_wishbone_tx_fifo_n1395, p_wishbone_tx_fifo_n1396, 
        p_wishbone_tx_fifo_n1397, p_wishbone_tx_fifo_n1398, 
        p_wishbone_tx_fifo_n1399, p_wishbone_tx_fifo_n1400, 
        p_wishbone_tx_fifo_n1401, p_wishbone_tx_fifo_n1402, 
        p_wishbone_tx_fifo_n1403, p_wishbone_tx_fifo_n1404, 
        p_wishbone_tx_fifo_n1405, p_wishbone_tx_fifo_n1406, 
        p_wishbone_tx_fifo_n1407, p_wishbone_tx_fifo_n1408, 
        p_wishbone_tx_fifo_n1409, p_wishbone_tx_fifo_n1410, 
        p_wishbone_tx_fifo_n1411, p_wishbone_tx_fifo_n1412, 
        p_wishbone_tx_fifo_n1413, p_wishbone_tx_fifo_n1414, 
        p_wishbone_tx_fifo_n1415, p_wishbone_tx_fifo_n1416, 
        p_wishbone_tx_fifo_n1417, p_wishbone_tx_fifo_n1418, 
        p_wishbone_tx_fifo_n1419, p_wishbone_tx_fifo_n1420, 
        p_wishbone_tx_fifo_n1421, p_wishbone_tx_fifo_n1422, 
        p_wishbone_tx_fifo_n1423, p_wishbone_tx_fifo_n1424, 
        p_wishbone_tx_fifo_n1425, p_wishbone_tx_fifo_n1426, 
        p_wishbone_tx_fifo_n1427, p_wishbone_tx_fifo_n1428, 
        p_wishbone_tx_fifo_n1429, p_wishbone_tx_fifo_n1430, 
        p_wishbone_tx_fifo_n1431, p_wishbone_tx_fifo_n1432, 
        p_wishbone_tx_fifo_n1433, p_wishbone_tx_fifo_n1434, 
        p_wishbone_tx_fifo_n1435, p_wishbone_tx_fifo_n1436, 
        p_wishbone_tx_fifo_n1437, p_wishbone_tx_fifo_n1438, 
        p_wishbone_tx_fifo_n1439, p_wishbone_tx_fifo_n1440, 
        p_wishbone_tx_fifo_n1441, p_wishbone_tx_fifo_n1442, 
        p_wishbone_tx_fifo_n1443, p_wishbone_tx_fifo_n1444, 
        p_wishbone_tx_fifo_n1445, p_wishbone_tx_fifo_n1446, 
        p_wishbone_tx_fifo_n1447, p_wishbone_tx_fifo_n1448, 
        p_wishbone_tx_fifo_n1449, p_wishbone_tx_fifo_n1450, 
        p_wishbone_tx_fifo_n1451, p_wishbone_tx_fifo_n1452, 
        p_wishbone_tx_fifo_n1453, p_wishbone_tx_fifo_n1454, 
        p_wishbone_tx_fifo_n1455, p_wishbone_tx_fifo_n1456, 
        p_wishbone_tx_fifo_n1457, p_wishbone_tx_fifo_n1458, 
        p_wishbone_tx_fifo_n1459, p_wishbone_tx_fifo_n1460, 
        p_wishbone_tx_fifo_n1461, p_wishbone_tx_fifo_n1462, 
        p_wishbone_tx_fifo_n1463, p_wishbone_tx_fifo_n1464, 
        p_wishbone_tx_fifo_n1465, p_wishbone_tx_fifo_n1466, 
        p_wishbone_tx_fifo_n1467, p_wishbone_tx_fifo_n1468, 
        p_wishbone_tx_fifo_n1469, p_wishbone_tx_fifo_n1470, 
        p_wishbone_tx_fifo_n1471, p_wishbone_tx_fifo_n1472, 
        p_wishbone_tx_fifo_n1473, p_wishbone_tx_fifo_n1474, 
        p_wishbone_tx_fifo_n1475, p_wishbone_tx_fifo_n1476, 
        p_wishbone_tx_fifo_n1477, p_wishbone_tx_fifo_n1478, 
        p_wishbone_tx_fifo_n1479, p_wishbone_tx_fifo_n1480, 
        p_wishbone_tx_fifo_n1481, p_wishbone_tx_fifo_n1482, 
        p_wishbone_tx_fifo_n1483, p_wishbone_tx_fifo_n1484, 
        p_wishbone_tx_fifo_n1485, p_wishbone_tx_fifo_n1486, 
        p_wishbone_tx_fifo_n1487, p_wishbone_tx_fifo_n1488, 
        p_wishbone_tx_fifo_n1489, p_wishbone_tx_fifo_n1490, 
        p_wishbone_tx_fifo_n1491, p_wishbone_tx_fifo_n1492, 
        p_wishbone_tx_fifo_n1493, p_wishbone_tx_fifo_n1494, 
        p_wishbone_tx_fifo_n1495, p_wishbone_tx_fifo_n1496, 
        p_wishbone_tx_fifo_n1497, p_wishbone_tx_fifo_n1498, 
        p_wishbone_tx_fifo_n1499, p_wishbone_tx_fifo_n1500, 
        p_wishbone_tx_fifo_n1501, p_wishbone_tx_fifo_n1502, 
        p_wishbone_tx_fifo_n1503, p_wishbone_tx_fifo_n1504, 
        p_wishbone_tx_fifo_n1505, p_wishbone_tx_fifo_n1506, 
        p_wishbone_tx_fifo_n1507, p_wishbone_tx_fifo_n1508, 
        p_wishbone_tx_fifo_n1509, p_wishbone_tx_fifo_n1510, 
        p_wishbone_tx_fifo_n1511, p_wishbone_tx_fifo_n1512, 
        p_wishbone_tx_fifo_n1513, p_wishbone_tx_fifo_n1514, 
        p_wishbone_tx_fifo_n1515, p_wishbone_tx_fifo_n1516, 
        p_wishbone_tx_fifo_n1517, p_wishbone_tx_fifo_n1518, 
        p_wishbone_tx_fifo_n1519, p_wishbone_tx_fifo_n1520, 
        p_wishbone_tx_fifo_n1521, p_wishbone_tx_fifo_n1522, 
        p_wishbone_tx_fifo_n1523, p_wishbone_tx_fifo_n1524, 
        p_wishbone_tx_fifo_n1525, p_wishbone_tx_fifo_n1526, 
        p_wishbone_tx_fifo_n1527, p_wishbone_tx_fifo_n1528, 
        p_wishbone_tx_fifo_n1529, p_wishbone_tx_fifo_n1530, 
        p_wishbone_tx_fifo_n1531, p_wishbone_tx_fifo_n1532, 
        p_wishbone_tx_fifo_n1533, p_wishbone_tx_fifo_n1534, 
        p_wishbone_tx_fifo_n1535, p_wishbone_tx_fifo_n1536, 
        p_wishbone_tx_fifo_n1537, p_wishbone_tx_fifo_n1538, 
        p_wishbone_tx_fifo_n1539, p_wishbone_tx_fifo_n1540, 
        p_wishbone_tx_fifo_n1541, p_wishbone_tx_fifo_n1542, 
        p_wishbone_tx_fifo_n1543, p_wishbone_tx_fifo_n1544, 
        p_wishbone_tx_fifo_n1545, p_wishbone_tx_fifo_n1546, 
        p_wishbone_tx_fifo_n1547, p_wishbone_tx_fifo_n1548, 
        p_wishbone_tx_fifo_n1549, p_wishbone_tx_fifo_n1550, 
        p_wishbone_tx_fifo_n1551, p_wishbone_tx_fifo_n1552, 
        p_wishbone_tx_fifo_n1553, p_wishbone_tx_fifo_n1554, 
        p_wishbone_tx_fifo_n1555, p_wishbone_tx_fifo_n1556, 
        p_wishbone_tx_fifo_n1557, p_wishbone_tx_fifo_n1558, 
        p_wishbone_tx_fifo_n1559, p_wishbone_tx_fifo_n1560, 
        p_wishbone_tx_fifo_n1561, p_wishbone_tx_fifo_n1562, 
        p_wishbone_tx_fifo_n1563, p_wishbone_tx_fifo_n1564, 
        p_wishbone_tx_fifo_n1565, p_wishbone_tx_fifo_n1566, 
        p_wishbone_tx_fifo_n1567, p_wishbone_tx_fifo_n1568, 
        p_wishbone_tx_fifo_n1569, p_wishbone_tx_fifo_n1570, 
        p_wishbone_tx_fifo_n1571, p_wishbone_tx_fifo_n1572, 
        p_wishbone_tx_fifo_n1573, p_wishbone_tx_fifo_n1574, 
        p_wishbone_tx_fifo_n1575, p_wishbone_tx_fifo_n1576, 
        p_wishbone_tx_fifo_n1577, p_wishbone_tx_fifo_n1578, 
        p_wishbone_tx_fifo_n1579, p_wishbone_tx_fifo_n1580, 
        p_wishbone_tx_fifo_n1581, p_wishbone_tx_fifo_n1582, 
        p_wishbone_tx_fifo_n1583, p_wishbone_tx_fifo_n1584, 
        p_wishbone_tx_fifo_n1585, p_wishbone_tx_fifo_n1586, 
        p_wishbone_tx_fifo_n1587, p_wishbone_tx_fifo_n1588, 
        p_wishbone_tx_fifo_n1589, p_wishbone_tx_fifo_n1590, 
        p_wishbone_tx_fifo_n1591, p_wishbone_tx_fifo_n1592, 
        p_wishbone_tx_fifo_n1593, p_wishbone_tx_fifo_n1594, 
        p_wishbone_tx_fifo_n1595, p_wishbone_tx_fifo_n1596, 
        p_wishbone_tx_fifo_n1597, p_wishbone_tx_fifo_n1598, 
        p_wishbone_tx_fifo_n1599, p_wishbone_tx_fifo_n1600, 
        p_wishbone_tx_fifo_n1601, p_wishbone_tx_fifo_n1602, 
        p_wishbone_tx_fifo_n1603, p_wishbone_tx_fifo_n1604, 
        p_wishbone_tx_fifo_n1605, p_wishbone_tx_fifo_n1606, 
        p_wishbone_tx_fifo_n1607, p_wishbone_tx_fifo_n1608, 
        p_wishbone_tx_fifo_n1609, p_wishbone_tx_fifo_n1610, 
        p_wishbone_tx_fifo_n1611, p_wishbone_tx_fifo_n1612, 
        p_wishbone_tx_fifo_n1613, p_wishbone_tx_fifo_n1614, 
        p_wishbone_tx_fifo_n1615, p_wishbone_tx_fifo_n1616, 
        p_wishbone_tx_fifo_n1617, p_wishbone_tx_fifo_n1618, 
        p_wishbone_tx_fifo_n1619, p_wishbone_tx_fifo_n1620, 
        p_wishbone_tx_fifo_n1621, p_wishbone_tx_fifo_n1622, 
        p_wishbone_tx_fifo_n1623, p_wishbone_tx_fifo_n1624, 
        p_wishbone_tx_fifo_n1625, p_wishbone_tx_fifo_n1626, 
        p_wishbone_tx_fifo_n1627, p_wishbone_tx_fifo_n1628, 
        p_wishbone_tx_fifo_n1629, p_wishbone_tx_fifo_n1630, 
        p_wishbone_tx_fifo_n1631, p_wishbone_tx_fifo_n1632, 
        p_wishbone_tx_fifo_n1633, p_wishbone_tx_fifo_n1634, 
        p_wishbone_tx_fifo_n1635, p_wishbone_tx_fifo_n1636, 
        p_wishbone_tx_fifo_n1637, p_wishbone_tx_fifo_n1638, 
        p_wishbone_tx_fifo_n1639, p_wishbone_tx_fifo_n1640, 
        p_wishbone_tx_fifo_n1641, p_wishbone_tx_fifo_n1642, 
        p_wishbone_tx_fifo_n1643, p_wishbone_tx_fifo_n1644, 
        p_wishbone_tx_fifo_n1645, p_wishbone_tx_fifo_n1646, 
        p_wishbone_tx_fifo_n1647, p_wishbone_tx_fifo_n1648, 
        p_wishbone_tx_fifo_n1649, p_wishbone_tx_fifo_n1650, 
        p_wishbone_tx_fifo_n1651, p_wishbone_tx_fifo_n1652, 
        p_wishbone_tx_fifo_n1653, p_wishbone_tx_fifo_n1654, 
        p_wishbone_tx_fifo_n1655, p_wishbone_tx_fifo_n1656, 
        p_wishbone_tx_fifo_n1657, p_wishbone_tx_fifo_n1658, 
        p_wishbone_tx_fifo_n1659, p_wishbone_tx_fifo_n1660, 
        p_wishbone_tx_fifo_n1661, p_wishbone_tx_fifo_n1662, 
        p_wishbone_tx_fifo_n1663, p_wishbone_tx_fifo_n1664, 
        p_wishbone_tx_fifo_n1665, p_wishbone_tx_fifo_n1666, 
        p_wishbone_tx_fifo_n1667, p_wishbone_tx_fifo_n1668, 
        p_wishbone_tx_fifo_n1669, p_wishbone_tx_fifo_n1670, 
        p_wishbone_tx_fifo_n1671, p_wishbone_tx_fifo_n1672, 
        p_wishbone_tx_fifo_n1673, p_wishbone_tx_fifo_n1674, 
        p_wishbone_tx_fifo_n1675, p_wishbone_tx_fifo_n1676, 
        p_wishbone_tx_fifo_n1677, p_wishbone_tx_fifo_n1678, 
        p_wishbone_tx_fifo_n1679, p_wishbone_tx_fifo_n1680, 
        p_wishbone_tx_fifo_n1681, p_wishbone_tx_fifo_n1682, 
        p_wishbone_tx_fifo_n1683, p_wishbone_tx_fifo_n1684, 
        p_wishbone_tx_fifo_n1685, p_wishbone_tx_fifo_n1686, 
        p_wishbone_tx_fifo_n1687, p_wishbone_tx_fifo_n1688, 
        p_wishbone_tx_fifo_n1689, p_wishbone_tx_fifo_n1690, 
        p_wishbone_tx_fifo_n1691, p_wishbone_tx_fifo_n1692, 
        p_wishbone_tx_fifo_n1693, p_wishbone_tx_fifo_n1694, 
        p_wishbone_tx_fifo_n1695, p_wishbone_tx_fifo_n1696, 
        p_wishbone_tx_fifo_n1697, p_wishbone_tx_fifo_n1698, 
        p_wishbone_tx_fifo_n1699, p_wishbone_tx_fifo_n1700, 
        p_wishbone_tx_fifo_n1701, p_wishbone_tx_fifo_n1702, 
        p_wishbone_tx_fifo_n1703, p_wishbone_tx_fifo_n1704, 
        p_wishbone_tx_fifo_n1705, p_wishbone_tx_fifo_n1706, 
        p_wishbone_tx_fifo_n1707, p_wishbone_tx_fifo_n1708, 
        p_wishbone_tx_fifo_n1709, p_wishbone_tx_fifo_n1710, 
        p_wishbone_tx_fifo_n1711, p_wishbone_tx_fifo_n1712, 
        p_wishbone_tx_fifo_n1713, p_wishbone_tx_fifo_n1714, 
        p_wishbone_tx_fifo_n1715, p_wishbone_tx_fifo_n1716, 
        p_wishbone_tx_fifo_n1717, p_wishbone_tx_fifo_n1718, 
        p_wishbone_tx_fifo_n1719, p_wishbone_tx_fifo_n1720, 
        p_wishbone_tx_fifo_n1721, p_wishbone_tx_fifo_n1722, 
        p_wishbone_tx_fifo_n1723, p_wishbone_tx_fifo_n1724, 
        p_wishbone_tx_fifo_n1725, p_wishbone_tx_fifo_n1726, 
        p_wishbone_tx_fifo_n1727, p_wishbone_tx_fifo_n1728, 
        p_wishbone_tx_fifo_n1729, p_wishbone_tx_fifo_n1730, 
        p_wishbone_tx_fifo_n1731, p_wishbone_tx_fifo_n1732, 
        p_wishbone_tx_fifo_n1733, p_wishbone_tx_fifo_n1734, 
        p_wishbone_tx_fifo_n1735, p_wishbone_tx_fifo_n1736, 
        p_wishbone_tx_fifo_n1737, p_wishbone_tx_fifo_n1738, 
        p_wishbone_tx_fifo_n1739, p_wishbone_tx_fifo_n1740, 
        p_wishbone_tx_fifo_n1741, p_wishbone_tx_fifo_n1742, 
        p_wishbone_tx_fifo_n1743, p_wishbone_tx_fifo_n1744, 
        p_wishbone_tx_fifo_n1745, p_wishbone_tx_fifo_n1746, 
        p_wishbone_tx_fifo_n1747, p_wishbone_tx_fifo_n1748, 
        p_wishbone_tx_fifo_n1749, p_wishbone_tx_fifo_n1750, 
        p_wishbone_tx_fifo_n1751, p_wishbone_tx_fifo_n1752, 
        p_wishbone_tx_fifo_n1753, n36050, n36051, n36052, n36053, n36054, 
        n36055, n36056, n36057, n36042, n36043, n36044, n36045, n36046, n36047, 
        n36048, n36049, n36034, n36035, n36036, n36037, n36038, n36039, n36040, 
        n36041, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, 
        n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36010, 
        n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36002, n36003, 
        n36004, n36005, n36006, n36007, n36008, n36009, n35994, n35995, n35996, 
        n35997, n35998, n35999, n36000, n36001, n35986, n35987, n35988, n35989, 
        n35990, n35991, n35992, n35993, n35978, n35979, n35980, n35981, n35982, 
        n35983, n35984, n35985, n35970, n35971, n35972, n35973, n35974, n35975, 
        n35976, n35977, n35962, n35963, n35964, n35965, n35966, n35967, n35968, 
        n35969, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, 
        n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35938, 
        n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35930, n35931, 
        n35932, n35933, n35934, n35935, n35936, n35937, n35922, n35923, n35924, 
        n35925, n35926, n35927, n35928, n35929, n35914, n35915, n35916, n35917, 
        n35918, n35919, n35920, n35921, n35906, n35907, n35908, n35909, n35910, 
        n35911, n35912, n35913, n35898, n35899, n35900, n35901, n35902, n35903, 
        n35904, n35905, n35897, n33925, n35892, n33930, n35893, n35894, n33926, 
        n35895, n35896, n35885, n35886, n35887, n35888, n35889, n35890, n35884, 
        n35891, n35883, n35882, n35877, n35878, n35879, n35880, n35881, 
        p_rxethmac1_crcrx_N25, p_rxethmac1_crcrx_N21, p_rxethmac1_crcrx_N17, 
        p_rxethmac1_crcrx_N13, p_rxethmac1_crcrx_N9, p_rxethmac1_crcrx_N5, 
        p_rxethmac1_crcrx_N8, p_rxethmac1_crcrx_N26, p_rxethmac1_crcrx_N22, 
        p_rxethmac1_crcrx_N18, p_rxethmac1_crcrx_N14, p_rxethmac1_crcrx_N10, 
        p_rxethmac1_crcrx_N6, p_rxethmac1_crcrx_N34, p_rxethmac1_crcrx_N30, 
        p_rxethmac1_crcrx_N4, p_rxethmac1_crcrx_N32, p_rxethmac1_crcrx_N28, 
        p_rxethmac1_crcrx_N24, p_rxethmac1_crcrx_N20, p_rxethmac1_crcrx_N16, 
        p_rxethmac1_crcrx_N12, p_rxethmac1_crcrx_N33, p_rxethmac1_crcrx_N29, 
        p_rxethmac1_crcrx_N31, p_rxethmac1_crcrx_N27, p_rxethmac1_crcrx_N23, 
        p_rxethmac1_crcrx_N19, p_rxethmac1_crcrx_N15, p_rxethmac1_crcrx_N11, 
        p_rxethmac1_crcrx_N7, p_rxethmac1_crcrx_N3, p_wishbone_rx_fifo_N623, 
        p_wishbone_rx_fifo_N624, p_wishbone_rx_fifo_N625, 
        p_wishbone_rx_fifo_N626, p_wishbone_rx_fifo_N627, 
        p_wishbone_rx_fifo_N628, p_wishbone_rx_fifo_N629, 
        p_wishbone_rx_fifo_N630, p_wishbone_rx_fifo_N631, 
        p_wishbone_rx_fifo_N632, p_wishbone_rx_fifo_N633, 
        p_wishbone_rx_fifo_N634, p_wishbone_rx_fifo_N635, 
        p_wishbone_rx_fifo_N636, p_wishbone_rx_fifo_N637, 
        p_wishbone_rx_fifo_N638, p_wishbone_rx_fifo_N639, 
        p_wishbone_rx_fifo_N640, p_wishbone_rx_fifo_N641, 
        p_wishbone_rx_fifo_N642, p_wishbone_rx_fifo_N643, 
        p_wishbone_rx_fifo_N644, p_wishbone_rx_fifo_N645, 
        p_wishbone_rx_fifo_N646, p_wishbone_rx_fifo_N647, 
        p_wishbone_rx_fifo_N648, p_wishbone_rx_fifo_N649, 
        p_wishbone_rx_fifo_N650, p_wishbone_rx_fifo_N651, 
        p_wishbone_rx_fifo_N652, p_wishbone_rx_fifo_N653, 
        p_wishbone_rx_fifo_N654, n33944, n33945, n33946, n33947, n33948, 
        n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, 
        n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, 
        n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, 
        n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, 
        n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, 
        n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, 
        n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, 
        n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, 
        n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, 
        n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, 
        n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, 
        n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, 
        n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, 
        n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, 
        n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, 
        n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, 
        n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, 
        n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, 
        n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, 
        n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, 
        n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, 
        n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, 
        n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, 
        n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, 
        n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, 
        n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, 
        n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, 
        n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, 
        n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, 
        n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, 
        n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, 
        n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, 
        n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, 
        n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, 
        n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, 
        n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, 
        n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, 
        n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, 
        n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, 
        n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, 
        n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, 
        n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, 
        n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, 
        n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, 
        n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, 
        n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, 
        n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, 
        n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, 
        n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, 
        n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, 
        n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, 
        n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, 
        n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, 
        n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, 
        n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, 
        n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, 
        n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, 
        n34462, n34463, n34464, n34465, n34466, n34467, n34468 );
  input wb_dat_i_0, wb_dat_i_1, wb_dat_i_2, wb_dat_i_3, wb_dat_i_4, wb_dat_i_5,
         wb_dat_i_6, wb_dat_i_7, wb_dat_i_8, wb_dat_i_9, wb_dat_i_10,
         wb_dat_i_11, wb_dat_i_12, wb_dat_i_13, wb_dat_i_14, wb_dat_i_15,
         wb_dat_i_16, wb_dat_i_17, wb_dat_i_18, wb_dat_i_19, wb_dat_i_20,
         wb_dat_i_21, wb_dat_i_22, wb_dat_i_23, wb_dat_i_24, wb_dat_i_25,
         wb_dat_i_26, wb_dat_i_27, wb_dat_i_28, wb_dat_i_29, wb_dat_i_30,
         wb_dat_i_31, wb_adr_i_2, wb_adr_i_3, wb_adr_i_4, wb_adr_i_5,
         wb_adr_i_6, wb_adr_i_7, wb_adr_i_8, wb_adr_i_9, wb_adr_i_10,
         wb_adr_i_11, wb_sel_i_0, wb_sel_i_1, wb_sel_i_2, wb_sel_i_3,
         m_wb_dat_i_0, m_wb_dat_i_1, m_wb_dat_i_2, m_wb_dat_i_3, m_wb_dat_i_4,
         m_wb_dat_i_5, m_wb_dat_i_6, m_wb_dat_i_7, m_wb_dat_i_8, m_wb_dat_i_9,
         m_wb_dat_i_10, m_wb_dat_i_11, m_wb_dat_i_12, m_wb_dat_i_13,
         m_wb_dat_i_14, m_wb_dat_i_15, m_wb_dat_i_16, m_wb_dat_i_17,
         m_wb_dat_i_18, m_wb_dat_i_19, m_wb_dat_i_20, m_wb_dat_i_21,
         m_wb_dat_i_22, m_wb_dat_i_23, m_wb_dat_i_24, m_wb_dat_i_25,
         m_wb_dat_i_26, m_wb_dat_i_27, m_wb_dat_i_28, m_wb_dat_i_29,
         m_wb_dat_i_30, m_wb_dat_i_31, mrxd_pad_i_0, mrxd_pad_i_1,
         mrxd_pad_i_2, mrxd_pad_i_3, wb_clk_i, wb_rst_i, wb_we_i, wb_cyc_i,
         wb_stb_i, m_wb_ack_i, m_wb_err_i, mtx_clk_pad_i, mrx_clk_pad_i,
         mrxdv_pad_i, mrxerr_pad_i, mcoll_pad_i, mcrs_pad_i, md_pad_i,
         BD_WB_DAT_O_0, BD_WB_DAT_O_1, BD_WB_DAT_O_2, BD_WB_DAT_O_3,
         BD_WB_DAT_O_4, BD_WB_DAT_O_5, BD_WB_DAT_O_6, BD_WB_DAT_O_7,
         BD_WB_DAT_O_8, BD_WB_DAT_O_9, BD_WB_DAT_O_10, BD_WB_DAT_O_11,
         BD_WB_DAT_O_12, BD_WB_DAT_O_13, BD_WB_DAT_O_14, BD_WB_DAT_O_15,
         BD_WB_DAT_O_16, BD_WB_DAT_O_17, BD_WB_DAT_O_18, BD_WB_DAT_O_19,
         BD_WB_DAT_O_20, BD_WB_DAT_O_21, BD_WB_DAT_O_22, BD_WB_DAT_O_23,
         BD_WB_DAT_O_24, BD_WB_DAT_O_25, BD_WB_DAT_O_26, BD_WB_DAT_O_27,
         BD_WB_DAT_O_28, BD_WB_DAT_O_29, BD_WB_DAT_O_30, BD_WB_DAT_O_31,
         CarrierSense_Tx1, CarrierSense_Tx2, Collision_Tx1, RxAbortRst,
         RxAbort_latch, RxAbort_sync1, RxAbort_wb, WillSendControlFrame_sync1,
         WillSendControlFrame_sync2, WillSendControlFrame_sync3, RstTxPauseRq,
         TxPauseRq_sync1, TxPauseRq_sync2, TxPauseRq_sync3, TPauseRq, RxEnSync,
         Collision_Tx2, WillTransmit_q, WillTransmit_q2, p_miim1_LatchByte_0,
         p_miim1_LatchByte0_d, p_miim1_LatchByte_1, p_miim1_LatchByte1_d,
         p_miim1_WriteOp, p_miim1_BitCounter_6, p_miim1_BitCounter_4,
         p_miim1_BitCounter_3, p_miim1_BitCounter_2, p_miim1_BitCounter_5,
         p_miim1_BitCounter_1, NValid_stat, UpdateMIIRX_DATAReg,
         p_miim1_WCtrlDataStart_q, p_miim1_RStatStart_q2,
         p_miim1_RStatStart_q1, RStatStart, p_miim1_WCtrlDataStart_q2,
         p_miim1_WCtrlDataStart_q1, WCtrlDataStart, p_miim1_EndBusy,
         p_miim1_InProgress_q3, p_miim1_InProgress_q2, p_miim1_InProgress_q1,
         p_miim1_InProgress, p_miim1_BitCounter_0, p_miim1_WCtrlData_q3,
         p_miim1_RStat_q3, p_miim1_SyncStatMdcEn, p_miim1_ScanStat_q2,
         p_ethreg1_INT_SOURCEOut_6, p_ethreg1_INT_SOURCEOut_5,
         p_ethreg1_INT_SOURCEOut_4, p_ethreg1_INT_SOURCEOut_3,
         p_ethreg1_INT_SOURCEOut_2, p_ethreg1_INT_SOURCEOut_1,
         p_ethreg1_INT_SOURCEOut_0, p_ethreg1_SetRxCIrq,
         p_ethreg1_ResetRxCIrq_sync2, p_ethreg1_SetRxCIrq_sync3,
         p_ethreg1_ResetRxCIrq_sync3, p_ethreg1_SetTxCIrq,
         p_ethreg1_SetTxCIrq_sync3, p_ethreg1_ResetTxCIrq_sync2,
         p_maccontrol1_MuxedDone, p_maccontrol1_MuxedAbort,
         p_maccontrol1_TxDoneInLatched, p_maccontrol1_TxAbortInLatched,
         p_maccontrol1_TxUsedDataOutDetected, RetryCnt_2, RetryCnt_1,
         p_txethmac1_PacketFinished, TxRetry, p_txethmac1_StatusLatch,
         p_txethmac1_ColWindow, p_txethmac1_StopExcessiveDeferOccured,
         TxUsedDataIn, RetryCnt_3, RetryCnt_0, p_txethmac1_PacketFinished_q,
         p_rxethmac1_Broadcast, p_rxethmac1_Multicast, RxEndFrm,
         p_rxethmac1_RxEndFrm_d, RxStartFrm, RxValid, RxData_7, RxData_6,
         RxData_5, RxData_4, RxData_3, RxData_2, RxData_1, RxData_0,
         p_rxethmac1_DelayData, p_rxethmac1_LatchedByte_0,
         p_rxethmac1_LatchedByte_1, p_rxethmac1_LatchedByte_2,
         p_rxethmac1_LatchedByte_3, p_rxethmac1_CrcHash_0,
         p_rxethmac1_CrcHash_1, p_rxethmac1_CrcHash_2, p_rxethmac1_CrcHash_3,
         p_rxethmac1_CrcHash_4, p_rxethmac1_CrcHash_5, p_rxethmac1_CrcHashGood,
         p_wishbone_Busy_IRQ_syncb1, p_wishbone_Busy_IRQ_sync3,
         p_wishbone_Busy_IRQ_syncb2, RxE_IRQ, RxB_IRQ, TxE_IRQ, TxB_IRQ,
         p_wishbone_RxStatusWriteLatched_syncb1,
         p_wishbone_RxStatusWriteLatched_syncb2, p_wishbone_RxPointerMSB_30,
         p_wishbone_RxPointerMSB_29, p_wishbone_RxPointerMSB_28,
         p_wishbone_RxPointerMSB_27, p_wishbone_RxPointerMSB_26,
         p_wishbone_RxPointerMSB_25, p_wishbone_RxPointerMSB_24,
         p_wishbone_RxPointerMSB_23, p_wishbone_RxPointerMSB_22,
         p_wishbone_RxPointerMSB_21, p_wishbone_RxPointerMSB_20,
         p_wishbone_RxPointerMSB_19, p_wishbone_RxPointerMSB_18,
         p_wishbone_RxPointerMSB_17, p_wishbone_RxPointerMSB_16,
         p_wishbone_RxPointerMSB_15, p_wishbone_RxPointerMSB_14,
         p_wishbone_RxPointerMSB_13, p_wishbone_RxPointerMSB_12,
         p_wishbone_RxPointerMSB_11, p_wishbone_RxPointerMSB_10,
         p_wishbone_RxPointerMSB_9, p_wishbone_RxPointerMSB_8,
         p_wishbone_RxPointerMSB_7, p_wishbone_RxPointerMSB_6,
         p_wishbone_RxPointerMSB_5, p_wishbone_RxPointerMSB_4,
         p_wishbone_RxPointerMSB_3, p_wishbone_RxPointerMSB_2,
         p_wishbone_RxPointerMSB_31, p_wishbone_TxPointerMSB_30,
         p_wishbone_TxPointerMSB_29, p_wishbone_TxPointerMSB_28,
         p_wishbone_TxPointerMSB_27, p_wishbone_TxPointerMSB_26,
         p_wishbone_TxPointerMSB_25, p_wishbone_TxPointerMSB_24,
         p_wishbone_TxPointerMSB_23, p_wishbone_TxPointerMSB_22,
         p_wishbone_TxPointerMSB_21, p_wishbone_TxPointerMSB_20,
         p_wishbone_TxPointerMSB_19, p_wishbone_TxPointerMSB_18,
         p_wishbone_TxPointerMSB_17, p_wishbone_TxPointerMSB_16,
         p_wishbone_TxPointerMSB_15, p_wishbone_TxPointerMSB_14,
         p_wishbone_TxPointerMSB_13, p_wishbone_TxPointerMSB_12,
         p_wishbone_TxPointerMSB_11, p_wishbone_TxPointerMSB_10,
         p_wishbone_TxPointerMSB_9, p_wishbone_TxPointerMSB_8,
         p_wishbone_TxPointerMSB_7, p_wishbone_TxPointerMSB_6,
         p_wishbone_TxPointerMSB_5, p_wishbone_TxPointerMSB_4,
         p_wishbone_TxPointerMSB_3, p_wishbone_TxPointerMSB_2,
         p_wishbone_TxPointerMSB_31, p_wishbone_BlockingIncrementTxPointer,
         p_wishbone_IncrTxPointer, p_wishbone_rx_burst_cnt_1,
         p_wishbone_rx_burst_cnt_0, p_wishbone_TxAbortPacketBlocked, TxData_7,
         p_wishbone_TxDataLatched_31, TxData_6, p_wishbone_TxDataLatched_30,
         TxData_5, p_wishbone_TxDataLatched_29, TxData_4,
         p_wishbone_TxDataLatched_28, TxData_3, p_wishbone_TxDataLatched_27,
         TxData_2, p_wishbone_TxDataLatched_26, TxData_1,
         p_wishbone_TxDataLatched_25, TxData_0, p_wishbone_TxDataLatched_24,
         p_wishbone_TxDataLatched_23, p_wishbone_TxDataLatched_22,
         p_wishbone_TxDataLatched_21, p_wishbone_TxDataLatched_20,
         p_wishbone_TxDataLatched_19, p_wishbone_TxDataLatched_18,
         p_wishbone_TxDataLatched_17, p_wishbone_TxDataLatched_16,
         p_wishbone_TxDataLatched_15, p_wishbone_TxDataLatched_14,
         p_wishbone_TxDataLatched_13, p_wishbone_TxDataLatched_12,
         p_wishbone_TxDataLatched_11, p_wishbone_TxDataLatched_10,
         p_wishbone_TxDataLatched_9, p_wishbone_TxDataLatched_8,
         p_wishbone_TxDataLatched_7, p_wishbone_TxDataLatched_6,
         p_wishbone_TxDataLatched_5, p_wishbone_TxDataLatched_4,
         p_wishbone_TxDataLatched_3, p_wishbone_TxDataLatched_2,
         p_wishbone_TxDataLatched_1, p_wishbone_TxDataLatched_0,
         p_wishbone_StartOccured, p_wishbone_TxByteCnt_1,
         p_wishbone_TxByteCnt_0, TxStartFrm, p_wishbone_TxStartFrm_syncb2,
         p_wishbone_TxEndFrm_wb, p_wishbone_ram_di_8, TxUnderRun,
         p_wishbone_TxUnderRun_sync1, p_wishbone_TxUnderRun_wb,
         p_wishbone_TxAbortPacket, p_wishbone_BlockingTxStatusWrite_sync3,
         p_wishbone_ram_addr_1, p_wishbone_ram_addr_7,
         p_wishbone_TxBDAddress_7, p_wishbone_ram_addr_6,
         p_wishbone_TxBDAddress_6, p_wishbone_ram_addr_5,
         p_wishbone_TxBDAddress_5, p_wishbone_ram_addr_4,
         p_wishbone_TxBDAddress_4, p_wishbone_ram_addr_3,
         p_wishbone_TxBDAddress_3, p_wishbone_ram_addr_2,
         p_wishbone_TxBDAddress_2, p_wishbone_TxBDAddress_1,
         p_wishbone_TxRetryPacket_NotCleared, p_wishbone_ram_addr_0,
         p_wishbone_TxPointerLSB_1, p_wishbone_TxPointerLSB_0,
         p_wishbone_ram_di_14, p_wishbone_ram_di_15, p_wishbone_ram_di_10,
         p_wishbone_ram_di_9, BDAck, p_wishbone_BDRead, p_wishbone_ram_di_31,
         p_wishbone_ram_di_30, p_wishbone_ram_di_29, p_wishbone_ram_di_28,
         p_wishbone_ram_di_27, p_wishbone_ram_di_26, p_wishbone_ram_di_25,
         p_wishbone_ram_di_24, p_wishbone_ram_di_23, p_wishbone_ram_di_22,
         p_wishbone_ram_di_21, p_wishbone_ram_di_20, p_wishbone_ram_di_19,
         p_wishbone_ram_di_18, p_wishbone_ram_di_17, p_wishbone_ram_di_16,
         p_wishbone_ram_di_13, p_wishbone_ram_di_12, p_wishbone_ram_di_11,
         p_wishbone_ram_di_7, p_wishbone_ram_di_5, p_wishbone_ram_di_4,
         p_wishbone_ram_di_3, p_wishbone_ram_di_2, p_wishbone_ram_di_1,
         p_wishbone_ram_di_0, p_wishbone_BDWrite_0, p_wishbone_BDWrite_1,
         p_wishbone_BDWrite_2, p_wishbone_BDWrite_3, p_wishbone_RxBDDataIn_14,
         p_wishbone_RxBDAddress_7, p_wishbone_RxBDAddress_6,
         p_wishbone_RxBDAddress_5, p_wishbone_RxBDAddress_4,
         p_wishbone_RxBDAddress_3, p_wishbone_RxBDAddress_2,
         p_wishbone_RxBDAddress_1, p_wishbone_RxBDDataIn_13,
         p_wishbone_ShiftEndedSync3, p_wishbone_RxDataLatched2_8,
         p_wishbone_RxDataLatched1_8, p_wishbone_RxDataLatched2_9,
         p_wishbone_RxDataLatched1_9, p_wishbone_RxDataLatched2_10,
         p_wishbone_RxDataLatched1_10, p_wishbone_RxDataLatched2_11,
         p_wishbone_RxDataLatched1_11, p_wishbone_RxDataLatched2_12,
         p_wishbone_RxDataLatched1_12, p_wishbone_RxDataLatched2_13,
         p_wishbone_RxDataLatched1_13, p_wishbone_RxDataLatched2_14,
         p_wishbone_RxDataLatched1_14, p_wishbone_RxDataLatched2_15,
         p_wishbone_RxDataLatched1_15, p_wishbone_RxDataLatched2_24,
         p_wishbone_RxDataLatched1_24, p_wishbone_RxDataLatched2_25,
         p_wishbone_RxDataLatched1_25, p_wishbone_RxDataLatched2_26,
         p_wishbone_RxDataLatched1_26, p_wishbone_RxDataLatched2_27,
         p_wishbone_RxDataLatched1_27, p_wishbone_RxDataLatched2_28,
         p_wishbone_RxDataLatched1_28, p_wishbone_RxDataLatched2_29,
         p_wishbone_RxDataLatched1_29, p_wishbone_RxDataLatched2_30,
         p_wishbone_RxDataLatched1_30, p_wishbone_RxDataLatched2_31,
         p_wishbone_RxDataLatched1_31, p_wishbone_RxDataLatched2_17,
         p_wishbone_RxDataLatched2_18, p_wishbone_RxDataLatched2_19,
         p_wishbone_RxDataLatched2_20, p_wishbone_RxDataLatched2_21,
         p_wishbone_RxDataLatched2_22, p_wishbone_RxDataLatched2_23,
         p_wishbone_RxDataLatched2_0, p_wishbone_RxDataLatched2_1,
         p_wishbone_RxDataLatched2_2, p_wishbone_RxDataLatched2_3,
         p_wishbone_RxDataLatched2_4, p_wishbone_RxDataLatched2_5,
         p_wishbone_RxDataLatched2_6, p_wishbone_RxDataLatched2_7,
         p_wishbone_WriteRxDataToFifoSync3, p_wishbone_RxByteCnt_1,
         p_wishbone_RxByteCnt_0, p_wishbone_ShiftWillEnd,
         p_wishbone_ShiftEndedSync_c2, p_wishbone_RxValidBytes_1,
         p_wishbone_RxValidBytes_0, p_wishbone_LastByteIn, p_wishbone_RxBDRead,
         p_wishbone_RxReady, p_wishbone_ShiftEnded,
         p_wishbone_RxDataLatched2_16, p_wishbone_RxDataLatched1_16,
         p_wishbone_RxDataLatched1_17, p_wishbone_RxDataLatched1_18,
         p_wishbone_RxDataLatched1_19, p_wishbone_RxDataLatched1_20,
         p_wishbone_RxDataLatched1_21, p_wishbone_RxDataLatched1_22,
         p_wishbone_RxDataLatched1_23, p_wishbone_RxPointerLSB_rst_0,
         p_wishbone_RxPointerLSB_rst_1, p_wishbone_RxPointerRead,
         p_wishbone_RxBDReady, p_wishbone_RxEn_q, p_wishbone_RxEn_needed,
         p_wishbone_WbEn_q, p_wishbone_LatchedTxLength_15,
         p_wishbone_LatchedTxLength_14, p_wishbone_LatchedTxLength_13,
         p_wishbone_LatchedTxLength_12, p_wishbone_LatchedTxLength_11,
         p_wishbone_LatchedTxLength_10, p_wishbone_LatchedTxLength_9,
         p_wishbone_LatchedTxLength_8, p_wishbone_LatchedTxLength_7,
         p_wishbone_LatchedTxLength_6, p_wishbone_LatchedTxLength_5,
         p_wishbone_LatchedTxLength_4, p_wishbone_LatchedTxLength_3,
         p_wishbone_LatchedTxLength_2, p_wishbone_LatchedTxLength_1,
         p_wishbone_LatchedTxLength_0, p_wishbone_BlockingTxBDRead,
         p_wishbone_TxBDReady, p_wishbone_ReadTxDataFromMemory,
         p_wishbone_TxLength_14, p_wishbone_TxLength_13,
         p_wishbone_TxLength_12, p_wishbone_TxLength_11,
         p_wishbone_TxLength_10, p_wishbone_TxLength_9, p_wishbone_TxLength_8,
         p_wishbone_TxLength_7, p_wishbone_TxLength_6, p_wishbone_TxLength_5,
         p_wishbone_TxLength_4, p_wishbone_TxLength_3, p_wishbone_TxLength_2,
         p_wishbone_TxValidBytesLatched_1, p_wishbone_TxLength_1,
         p_wishbone_TxLength_0, PerPacketCrcEn, PerPacketPad,
         p_wishbone_TxStatus_13, p_wishbone_TxStatus_14,
         p_wishbone_TxDonePacket_NotCleared, p_wishbone_TxEn_q,
         p_wishbone_TxEn_needed, p_wishbone_U3_U3_Z_0,
         p_wishbone_TxPointerLSB_rst_1, p_wishbone_TxPointerRead,
         p_wishbone_TxBDRead, p_wishbone_TxAbortPacket_NotCleared,
         p_wishbone_TxRetryPacketBlocked, p_wishbone_TxRetryPacket,
         p_wishbone_TxDonePacketBlocked, p_wishbone_TxDonePacket,
         p_wishbone_tx_burst_en, p_wishbone_tx_burst_cnt_2,
         p_wishbone_tx_burst_cnt_1, p_wishbone_tx_burst_cnt_0,
         p_wishbone_cyc_cleared, p_wishbone_MasterWbTX, p_wishbone_MasterWbRX,
         p_wishbone_rx_burst_en, p_wishbone_rx_burst_cnt_2,
         p_wishbone_BlockReadTxDataFromMemory,
         p_wishbone_ReadTxDataFromFifo_sync3,
         p_wishbone_ReadTxDataFromFifo_syncb3, p_wishbone_LastWord, TxEndFrm,
         p_wishbone_TxValidBytesLatched_0, p_wishbone_LatchValidBytes_q,
         p_wishbone_TxLength_15, p_wishbone_ram_di_6, p_wishbone_RxBDDataIn_6,
         p_wishbone_RxStatusIn_6, p_wishbone_RxBDDataIn_0,
         p_wishbone_RxBDDataIn_1, p_wishbone_RxBDDataIn_2,
         p_wishbone_RxBDDataIn_3, p_wishbone_RxBDDataIn_4,
         p_wishbone_RxBDDataIn_5, p_wishbone_RxBDDataIn_7,
         p_wishbone_RxBDDataIn_8, p_wishbone_RxBDDataIn_16,
         p_wishbone_RxBDDataIn_17, p_wishbone_RxBDDataIn_18,
         p_wishbone_RxBDDataIn_19, p_wishbone_RxBDDataIn_20,
         p_wishbone_RxBDDataIn_21, p_wishbone_RxBDDataIn_22,
         p_wishbone_RxBDDataIn_23, p_wishbone_RxBDDataIn_24,
         p_wishbone_RxBDDataIn_25, p_wishbone_RxBDDataIn_26,
         p_wishbone_RxBDDataIn_27, p_wishbone_RxBDDataIn_28,
         p_wishbone_RxBDDataIn_29, p_wishbone_RxBDDataIn_30,
         p_wishbone_RxBDDataIn_31, p_wishbone_RxAbortSyncb2,
         p_wishbone_RxAbortSync4, p_wishbone_RxEnableWindow,
         p_wishbone_SyncRxStartFrm_q2, p_wishbone_SyncRxStartFrm,
         p_wishbone_TxAbort_wb_q, p_wishbone_TxDone_wb_q,
         p_wishbone_TxRetry_wb_q, p_wishbone_TxAbort_q,
         p_wishbone_TxUsedData_q, p_wishbone_Flop, p_wishbone_TxRetry_q,
         p_wishbone_r_RxEn_q, p_wishbone_r_TxEn_q, CarrierSenseLost,
         DeferLatched, LateCollLatched, RetryLimit, RetryCntLatched_0,
         RetryCntLatched_1, RetryCntLatched_2, RetryCntLatched_3,
         ReceivedPacketTooBig, DribbleNibble, ShortFrame, RxLateCollision,
         p_macstatus1_RxColWindow, InvalidSymbol, ReceiveEnd, LatchedMRxErr,
         LatchedCrcError, p_miim1_clkgen_Counter_6, p_miim1_clkgen_Counter_5,
         p_miim1_clkgen_Counter_4, p_miim1_clkgen_Counter_3,
         p_miim1_clkgen_Counter_2, p_miim1_clkgen_Counter_1,
         p_miim1_clkgen_Counter_0, LinkFail, Prsd_0, Prsd_1, Prsd_2, Prsd_3,
         Prsd_4, Prsd_5, Prsd_6, Prsd_7, Prsd_8, Prsd_9, Prsd_10, Prsd_11,
         Prsd_12, Prsd_13, Prsd_14, Prsd_15, p_miim1_ShiftedBit,
         p_miim1_shftrg_ShiftReg_6, p_miim1_shftrg_ShiftReg_5,
         p_miim1_shftrg_ShiftReg_4, p_miim1_shftrg_ShiftReg_3,
         p_miim1_shftrg_ShiftReg_2, p_miim1_shftrg_ShiftReg_1,
         p_miim1_shftrg_ShiftReg_0, p_miim1_outctrl_Mdo_d,
         p_miim1_outctrl_Mdo_2d, p_miim1_outctrl_MdoEn_d,
         p_miim1_outctrl_MdoEn_2d, p_ethreg1_MODEROut_0, p_ethreg1_MODEROut_1,
         p_ethreg1_r_NoPre, r_Bro, p_ethreg1_r_Iam, r_Pro, r_IFG, r_LoopBck,
         r_NoBckof, r_ExDfrEn, r_FullD, p_ethreg1_MODEROut_11, r_DlyCrcEn,
         r_CrcEn, r_HugEn, r_Pad, r_RecSmall, p_ethreg1_INT_MASKOut_0,
         p_ethreg1_INT_MASKOut_1, p_ethreg1_INT_MASKOut_2,
         p_ethreg1_INT_MASKOut_3, p_ethreg1_INT_MASKOut_4,
         p_ethreg1_INT_MASKOut_5, p_ethreg1_INT_MASKOut_6, r_IPGT_0, r_IPGT_1,
         r_IPGT_2, r_IPGT_3, r_IPGT_4, r_IPGT_5, r_IPGT_6, r_IPGR1_0,
         r_IPGR1_1, r_IPGR1_2, r_IPGR1_3, r_IPGR1_4, r_IPGR1_5, r_IPGR1_6,
         r_MaxFL_8, r_MaxFL_9, r_MaxFL_10, r_MaxFL_11, r_MaxFL_12, r_MaxFL_13,
         r_MaxFL_14, r_MaxFL_15, p_txethmac1_txcounters1_N41,
         p_txethmac1_txcounters1_N42, r_MinFL_2, r_MinFL_3, r_MinFL_4,
         r_MinFL_5, r_MinFL_6, r_MinFL_7, r_CollValid_0, r_CollValid_1,
         r_CollValid_2, r_CollValid_3, r_CollValid_4, r_CollValid_5,
         r_MaxRet_0, r_MaxRet_1, r_MaxRet_2, r_MaxRet_3, r_PassAll, r_RxFlow,
         r_TxFlow, r_ClkDiv_0, r_ClkDiv_1, r_ClkDiv_2, r_ClkDiv_3, r_ClkDiv_4,
         r_ClkDiv_5, r_ClkDiv_6, r_ClkDiv_7, r_FIAD_0, r_FIAD_1, r_FIAD_2,
         r_FIAD_3, r_FIAD_4, p_ethreg1_MIIRX_DATAOut_0,
         p_ethreg1_MIIRX_DATAOut_1, p_ethreg1_MIIRX_DATAOut_2,
         p_ethreg1_MIIRX_DATAOut_3, p_ethreg1_MIIRX_DATAOut_4,
         p_ethreg1_MIIRX_DATAOut_5, p_ethreg1_MIIRX_DATAOut_6,
         p_ethreg1_MIIRX_DATAOut_7, p_ethreg1_MIIRX_DATAOut_8,
         p_ethreg1_MIIRX_DATAOut_9, p_ethreg1_MIIRX_DATAOut_10,
         p_ethreg1_MIIRX_DATAOut_11, p_ethreg1_MIIRX_DATAOut_12,
         p_ethreg1_MIIRX_DATAOut_13, p_ethreg1_MIIRX_DATAOut_14,
         p_ethreg1_MIIRX_DATAOut_15, ReceivedPauseFrm,
         p_maccontrol1_receivecontrol1_SlotTimer_4,
         p_maccontrol1_receivecontrol1_SlotTimer_3,
         p_maccontrol1_receivecontrol1_SlotTimer_2,
         p_maccontrol1_receivecontrol1_SlotTimer_1,
         p_maccontrol1_receivecontrol1_SlotTimer_5, p_maccontrol1_Pause,
         p_maccontrol1_receivecontrol1_PauseTimerEq0_sync2,
         p_maccontrol1_receivecontrol1_Divider2,
         p_maccontrol1_receivecontrol1_PauseTimer_15,
         p_maccontrol1_receivecontrol1_PauseTimer_14,
         p_maccontrol1_receivecontrol1_PauseTimer_13,
         p_maccontrol1_receivecontrol1_PauseTimer_12,
         p_maccontrol1_receivecontrol1_PauseTimer_11,
         p_maccontrol1_receivecontrol1_PauseTimer_10,
         p_maccontrol1_receivecontrol1_PauseTimer_9,
         p_maccontrol1_receivecontrol1_PauseTimer_8,
         p_maccontrol1_receivecontrol1_PauseTimer_7,
         p_maccontrol1_receivecontrol1_PauseTimer_6,
         p_maccontrol1_receivecontrol1_PauseTimer_5,
         p_maccontrol1_receivecontrol1_PauseTimer_4,
         p_maccontrol1_receivecontrol1_PauseTimer_3,
         p_maccontrol1_receivecontrol1_PauseTimer_2,
         p_maccontrol1_receivecontrol1_PauseTimer_1,
         p_maccontrol1_receivecontrol1_PauseTimer_0,
         p_maccontrol1_receivecontrol1_SlotTimer_0,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_0,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_1,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_2,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_3,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_4,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_5,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_6,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_7,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_8,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_9,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_10,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_11,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_12,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_13,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_14,
         p_maccontrol1_receivecontrol1_LatchedTimerValue_15,
         p_maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr,
         ControlFrmAddressOK, p_maccontrol1_receivecontrol1_OpCodeOK,
         p_maccontrol1_receivecontrol1_TypeLengthOK,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_0,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_1,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_2,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_3,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_4,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_5,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_6,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_7,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_8,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_9,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_10,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_11,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_12,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_13,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_14,
         p_maccontrol1_receivecontrol1_AssembledTimerValue_15,
         p_maccontrol1_receivecontrol1_ByteCnt_3,
         p_maccontrol1_receivecontrol1_ByteCnt_2,
         p_maccontrol1_receivecontrol1_ByteCnt_1,
         p_maccontrol1_receivecontrol1_ByteCnt_4,
         p_maccontrol1_receivecontrol1_DetectionWindow,
         p_maccontrol1_receivecontrol1_ByteCnt_0,
         p_maccontrol1_receivecontrol1_DlyCrcCnt_1,
         p_maccontrol1_receivecontrol1_DlyCrcCnt_2,
         p_maccontrol1_receivecontrol1_DlyCrcCnt_0,
         p_maccontrol1_ControlData_0, p_maccontrol1_ControlData_1,
         p_maccontrol1_ControlData_2, p_maccontrol1_ControlData_3,
         p_maccontrol1_ControlData_4, p_maccontrol1_ControlData_5,
         p_maccontrol1_ControlData_6, p_maccontrol1_ControlData_7,
         p_maccontrol1_transmitcontrol1_ByteCnt_4,
         p_maccontrol1_transmitcontrol1_ByteCnt_3,
         p_maccontrol1_transmitcontrol1_ByteCnt_2,
         p_maccontrol1_transmitcontrol1_ByteCnt_1,
         p_maccontrol1_transmitcontrol1_ByteCnt_5,
         p_maccontrol1_transmitcontrol1_DlyCrcCnt_2,
         p_maccontrol1_transmitcontrol1_DlyCrcCnt_1,
         p_maccontrol1_transmitcontrol1_DlyCrcCnt_0, p_maccontrol1_BlockTxDone,
         p_maccontrol1_SendingCtrlFrm,
         p_maccontrol1_transmitcontrol1_TxCtrlStartFrm_q,
         p_maccontrol1_CtrlMux, TxCtrlEndFrm,
         p_maccontrol1_transmitcontrol1_ControlEnd_q,
         p_maccontrol1_transmitcontrol1_ByteCnt_0,
         p_maccontrol1_transmitcontrol1_TxUsedDataIn_q,
         p_txethmac1_DlyCrcCnt_1, p_txethmac1_DlyCrcCnt_2,
         p_txethmac1_DlyCrcCnt_0, p_txethmac1_txcounters1_ByteCnt_14,
         p_txethmac1_txcounters1_ByteCnt_13,
         p_txethmac1_txcounters1_ByteCnt_12,
         p_txethmac1_txcounters1_ByteCnt_11,
         p_txethmac1_txcounters1_ByteCnt_10, p_txethmac1_ByteCnt_9,
         p_txethmac1_ByteCnt_8, p_txethmac1_ByteCnt_7, p_txethmac1_ByteCnt_6,
         p_txethmac1_ByteCnt_5, p_txethmac1_ByteCnt_4, p_txethmac1_ByteCnt_3,
         p_txethmac1_ByteCnt_2, p_txethmac1_ByteCnt_1,
         p_txethmac1_txcounters1_ByteCnt_15, p_txethmac1_ByteCnt_0,
         p_txethmac1_NibCnt_15, p_txethmac1_NibCnt_14, p_txethmac1_NibCnt_13,
         p_txethmac1_NibCnt_12, p_txethmac1_NibCnt_11, p_txethmac1_NibCnt_10,
         p_txethmac1_NibCnt_9, p_txethmac1_NibCnt_8, p_txethmac1_NibCnt_7,
         p_txethmac1_NibCnt_6, p_txethmac1_NibCnt_5, p_txethmac1_NibCnt_4,
         p_txethmac1_NibCnt_2, p_txethmac1_NibCnt_1, p_txethmac1_NibCnt_3,
         p_txethmac1_NibCnt_0, p_txethmac1_StateBackOff,
         p_txethmac1_StateJam_q, p_txethmac1_StatePAD, StateData_1,
         StateData_0, StatePreamble, p_txethmac1_StateFCS,
         p_txethmac1_StateIdle, p_txethmac1_StateDefer, p_txethmac1_StateIPG,
         p_txethmac1_txstatem1_Rule1, p_txethmac1_txcrc_Crc_22,
         p_txethmac1_txcrc_Crc_18, p_txethmac1_txcrc_Crc_14,
         p_txethmac1_txcrc_Crc_10, p_txethmac1_txcrc_Crc_6,
         p_txethmac1_txcrc_Crc_2, p_txethmac1_txcrc_Crc_5,
         p_txethmac1_txcrc_Crc_23, p_txethmac1_txcrc_Crc_19,
         p_txethmac1_txcrc_Crc_15, p_txethmac1_txcrc_Crc_11,
         p_txethmac1_txcrc_Crc_7, p_txethmac1_txcrc_Crc_3, p_txethmac1_Crc_31,
         p_txethmac1_txcrc_Crc_27, p_txethmac1_txcrc_Crc_1, p_txethmac1_Crc_29,
         p_txethmac1_txcrc_Crc_25, p_txethmac1_txcrc_Crc_21,
         p_txethmac1_txcrc_Crc_17, p_txethmac1_txcrc_Crc_13,
         p_txethmac1_txcrc_Crc_9, p_txethmac1_Crc_30, p_txethmac1_txcrc_Crc_26,
         p_txethmac1_Crc_28, p_txethmac1_txcrc_Crc_24,
         p_txethmac1_txcrc_Crc_20, p_txethmac1_txcrc_Crc_16,
         p_txethmac1_txcrc_Crc_12, p_txethmac1_txcrc_Crc_8,
         p_txethmac1_txcrc_Crc_4, p_txethmac1_txcrc_Crc_0,
         p_txethmac1_random1_RandomLatched_0,
         p_txethmac1_random1_RandomLatched_1,
         p_txethmac1_random1_RandomLatched_2,
         p_txethmac1_random1_RandomLatched_3,
         p_txethmac1_random1_RandomLatched_4,
         p_txethmac1_random1_RandomLatched_5,
         p_txethmac1_random1_RandomLatched_6,
         p_txethmac1_random1_RandomLatched_7,
         p_txethmac1_random1_RandomLatched_8,
         p_txethmac1_random1_RandomLatched_9, p_txethmac1_random1_x_9,
         RxStateSFD, RxStateData_1, RxStatePreamble, RxStateIdle,
         p_rxethmac1_StateDrop, p_rxethmac1_rxcounters1_ByteCnt_14,
         p_rxethmac1_rxcounters1_ByteCnt_13,
         p_rxethmac1_rxcounters1_ByteCnt_12,
         p_rxethmac1_rxcounters1_ByteCnt_11,
         p_rxethmac1_rxcounters1_ByteCnt_10, p_rxethmac1_rxcounters1_ByteCnt_9,
         p_rxethmac1_rxcounters1_ByteCnt_8, p_rxethmac1_rxcounters1_ByteCnt_7,
         p_rxethmac1_rxcounters1_ByteCnt_6, p_rxethmac1_rxcounters1_ByteCnt_5,
         p_rxethmac1_rxcounters1_ByteCnt_4, p_rxethmac1_rxcounters1_ByteCnt_3,
         p_rxethmac1_rxcounters1_ByteCnt_2, RxByteCnt_1,
         p_rxethmac1_rxcounters1_ByteCnt_15, RxByteCnt_0,
         p_rxethmac1_DlyCrcCnt_2, p_rxethmac1_DlyCrcCnt_1,
         p_rxethmac1_DlyCrcCnt_3, p_rxethmac1_DlyCrcCnt_0,
         p_rxethmac1_rxcounters1_IFGCounter_3,
         p_rxethmac1_rxcounters1_IFGCounter_2,
         p_rxethmac1_rxcounters1_IFGCounter_1,
         p_rxethmac1_rxcounters1_IFGCounter_4,
         p_rxethmac1_rxcounters1_IFGCounter_0, AddressMiss,
         p_rxethmac1_rxaddrcheck1_MulticastOK, RxAbort,
         p_rxethmac1_rxaddrcheck1_UnicastOK, p_wishbone_bd_ram_mem2_0_16,
         p_wishbone_bd_ram_mem2_0_17, p_wishbone_bd_ram_mem2_0_18,
         p_wishbone_bd_ram_mem2_0_19, p_wishbone_bd_ram_mem2_0_20,
         p_wishbone_bd_ram_mem2_0_21, p_wishbone_bd_ram_mem2_0_22,
         p_wishbone_bd_ram_mem2_0_23, p_wishbone_bd_ram_mem2_1_16,
         p_wishbone_bd_ram_mem2_1_17, p_wishbone_bd_ram_mem2_1_18,
         p_wishbone_bd_ram_mem2_1_19, p_wishbone_bd_ram_mem2_1_20,
         p_wishbone_bd_ram_mem2_1_21, p_wishbone_bd_ram_mem2_1_22,
         p_wishbone_bd_ram_mem2_1_23, p_wishbone_bd_ram_mem2_2_16,
         p_wishbone_bd_ram_mem2_2_17, p_wishbone_bd_ram_mem2_2_18,
         p_wishbone_bd_ram_mem2_2_19, p_wishbone_bd_ram_mem2_2_20,
         p_wishbone_bd_ram_mem2_2_21, p_wishbone_bd_ram_mem2_2_22,
         p_wishbone_bd_ram_mem2_2_23, p_wishbone_bd_ram_mem2_3_16,
         p_wishbone_bd_ram_mem2_3_17, p_wishbone_bd_ram_mem2_3_18,
         p_wishbone_bd_ram_mem2_3_19, p_wishbone_bd_ram_mem2_3_20,
         p_wishbone_bd_ram_mem2_3_21, p_wishbone_bd_ram_mem2_3_22,
         p_wishbone_bd_ram_mem2_3_23, p_wishbone_bd_ram_mem2_4_16,
         p_wishbone_bd_ram_mem2_4_17, p_wishbone_bd_ram_mem2_4_18,
         p_wishbone_bd_ram_mem2_4_19, p_wishbone_bd_ram_mem2_4_20,
         p_wishbone_bd_ram_mem2_4_21, p_wishbone_bd_ram_mem2_4_22,
         p_wishbone_bd_ram_mem2_4_23, p_wishbone_bd_ram_mem2_5_16,
         p_wishbone_bd_ram_mem2_5_17, p_wishbone_bd_ram_mem2_5_18,
         p_wishbone_bd_ram_mem2_5_19, p_wishbone_bd_ram_mem2_5_20,
         p_wishbone_bd_ram_mem2_5_21, p_wishbone_bd_ram_mem2_5_22,
         p_wishbone_bd_ram_mem2_5_23, p_wishbone_bd_ram_mem2_6_16,
         p_wishbone_bd_ram_mem2_6_17, p_wishbone_bd_ram_mem2_6_18,
         p_wishbone_bd_ram_mem2_6_19, p_wishbone_bd_ram_mem2_6_20,
         p_wishbone_bd_ram_mem2_6_21, p_wishbone_bd_ram_mem2_6_22,
         p_wishbone_bd_ram_mem2_6_23, p_wishbone_bd_ram_mem2_7_16,
         p_wishbone_bd_ram_mem2_7_17, p_wishbone_bd_ram_mem2_7_18,
         p_wishbone_bd_ram_mem2_7_19, p_wishbone_bd_ram_mem2_7_20,
         p_wishbone_bd_ram_mem2_7_21, p_wishbone_bd_ram_mem2_7_22,
         p_wishbone_bd_ram_mem2_7_23, p_wishbone_bd_ram_mem2_8_16,
         p_wishbone_bd_ram_mem2_8_17, p_wishbone_bd_ram_mem2_8_18,
         p_wishbone_bd_ram_mem2_8_19, p_wishbone_bd_ram_mem2_8_20,
         p_wishbone_bd_ram_mem2_8_21, p_wishbone_bd_ram_mem2_8_22,
         p_wishbone_bd_ram_mem2_8_23, p_wishbone_bd_ram_mem2_9_16,
         p_wishbone_bd_ram_mem2_9_17, p_wishbone_bd_ram_mem2_9_18,
         p_wishbone_bd_ram_mem2_9_19, p_wishbone_bd_ram_mem2_9_20,
         p_wishbone_bd_ram_mem2_9_21, p_wishbone_bd_ram_mem2_9_22,
         p_wishbone_bd_ram_mem2_9_23, p_wishbone_bd_ram_mem2_10_16,
         p_wishbone_bd_ram_mem2_10_17, p_wishbone_bd_ram_mem2_10_18,
         p_wishbone_bd_ram_mem2_10_19, p_wishbone_bd_ram_mem2_10_20,
         p_wishbone_bd_ram_mem2_10_21, p_wishbone_bd_ram_mem2_10_22,
         p_wishbone_bd_ram_mem2_10_23, p_wishbone_bd_ram_mem2_11_16,
         p_wishbone_bd_ram_mem2_11_17, p_wishbone_bd_ram_mem2_11_18,
         p_wishbone_bd_ram_mem2_11_19, p_wishbone_bd_ram_mem2_11_20,
         p_wishbone_bd_ram_mem2_11_21, p_wishbone_bd_ram_mem2_11_22,
         p_wishbone_bd_ram_mem2_11_23, p_wishbone_bd_ram_mem2_12_16,
         p_wishbone_bd_ram_mem2_12_17, p_wishbone_bd_ram_mem2_12_18,
         p_wishbone_bd_ram_mem2_12_19, p_wishbone_bd_ram_mem2_12_20,
         p_wishbone_bd_ram_mem2_12_21, p_wishbone_bd_ram_mem2_12_22,
         p_wishbone_bd_ram_mem2_12_23, p_wishbone_bd_ram_mem2_13_16,
         p_wishbone_bd_ram_mem2_13_17, p_wishbone_bd_ram_mem2_13_18,
         p_wishbone_bd_ram_mem2_13_19, p_wishbone_bd_ram_mem2_13_20,
         p_wishbone_bd_ram_mem2_13_21, p_wishbone_bd_ram_mem2_13_22,
         p_wishbone_bd_ram_mem2_13_23, p_wishbone_bd_ram_mem2_14_16,
         p_wishbone_bd_ram_mem2_14_17, p_wishbone_bd_ram_mem2_14_18,
         p_wishbone_bd_ram_mem2_14_19, p_wishbone_bd_ram_mem2_14_20,
         p_wishbone_bd_ram_mem2_14_21, p_wishbone_bd_ram_mem2_14_22,
         p_wishbone_bd_ram_mem2_14_23, p_wishbone_bd_ram_mem2_15_16,
         p_wishbone_bd_ram_mem2_15_17, p_wishbone_bd_ram_mem2_15_18,
         p_wishbone_bd_ram_mem2_15_19, p_wishbone_bd_ram_mem2_15_20,
         p_wishbone_bd_ram_mem2_15_21, p_wishbone_bd_ram_mem2_15_22,
         p_wishbone_bd_ram_mem2_15_23, p_wishbone_bd_ram_mem2_16_16,
         p_wishbone_bd_ram_mem2_16_17, p_wishbone_bd_ram_mem2_16_18,
         p_wishbone_bd_ram_mem2_16_19, p_wishbone_bd_ram_mem2_16_20,
         p_wishbone_bd_ram_mem2_16_21, p_wishbone_bd_ram_mem2_16_22,
         p_wishbone_bd_ram_mem2_16_23, p_wishbone_bd_ram_mem2_17_16,
         p_wishbone_bd_ram_mem2_17_17, p_wishbone_bd_ram_mem2_17_18,
         p_wishbone_bd_ram_mem2_17_19, p_wishbone_bd_ram_mem2_17_20,
         p_wishbone_bd_ram_mem2_17_21, p_wishbone_bd_ram_mem2_17_22,
         p_wishbone_bd_ram_mem2_17_23, p_wishbone_bd_ram_mem2_18_16,
         p_wishbone_bd_ram_mem2_18_17, p_wishbone_bd_ram_mem2_18_18,
         p_wishbone_bd_ram_mem2_18_19, p_wishbone_bd_ram_mem2_18_20,
         p_wishbone_bd_ram_mem2_18_21, p_wishbone_bd_ram_mem2_18_22,
         p_wishbone_bd_ram_mem2_18_23, p_wishbone_bd_ram_mem2_19_16,
         p_wishbone_bd_ram_mem2_19_17, p_wishbone_bd_ram_mem2_19_18,
         p_wishbone_bd_ram_mem2_19_19, p_wishbone_bd_ram_mem2_19_20,
         p_wishbone_bd_ram_mem2_19_21, p_wishbone_bd_ram_mem2_19_22,
         p_wishbone_bd_ram_mem2_19_23, p_wishbone_bd_ram_mem2_20_16,
         p_wishbone_bd_ram_mem2_20_17, p_wishbone_bd_ram_mem2_20_18,
         p_wishbone_bd_ram_mem2_20_19, p_wishbone_bd_ram_mem2_20_20,
         p_wishbone_bd_ram_mem2_20_21, p_wishbone_bd_ram_mem2_20_22,
         p_wishbone_bd_ram_mem2_20_23, p_wishbone_bd_ram_mem2_21_16,
         p_wishbone_bd_ram_mem2_21_17, p_wishbone_bd_ram_mem2_21_18,
         p_wishbone_bd_ram_mem2_21_19, p_wishbone_bd_ram_mem2_21_20,
         p_wishbone_bd_ram_mem2_21_21, p_wishbone_bd_ram_mem2_21_22,
         p_wishbone_bd_ram_mem2_21_23, p_wishbone_bd_ram_mem2_22_16,
         p_wishbone_bd_ram_mem2_22_17, p_wishbone_bd_ram_mem2_22_18,
         p_wishbone_bd_ram_mem2_22_19, p_wishbone_bd_ram_mem2_22_20,
         p_wishbone_bd_ram_mem2_22_21, p_wishbone_bd_ram_mem2_22_22,
         p_wishbone_bd_ram_mem2_22_23, p_wishbone_bd_ram_mem2_23_16,
         p_wishbone_bd_ram_mem2_23_17, p_wishbone_bd_ram_mem2_23_18,
         p_wishbone_bd_ram_mem2_23_19, p_wishbone_bd_ram_mem2_23_20,
         p_wishbone_bd_ram_mem2_23_21, p_wishbone_bd_ram_mem2_23_22,
         p_wishbone_bd_ram_mem2_23_23, p_wishbone_bd_ram_mem2_24_16,
         p_wishbone_bd_ram_mem2_24_17, p_wishbone_bd_ram_mem2_24_18,
         p_wishbone_bd_ram_mem2_24_19, p_wishbone_bd_ram_mem2_24_20,
         p_wishbone_bd_ram_mem2_24_21, p_wishbone_bd_ram_mem2_24_22,
         p_wishbone_bd_ram_mem2_24_23, p_wishbone_bd_ram_mem2_25_16,
         p_wishbone_bd_ram_mem2_25_17, p_wishbone_bd_ram_mem2_25_18,
         p_wishbone_bd_ram_mem2_25_19, p_wishbone_bd_ram_mem2_25_20,
         p_wishbone_bd_ram_mem2_25_21, p_wishbone_bd_ram_mem2_25_22,
         p_wishbone_bd_ram_mem2_25_23, p_wishbone_bd_ram_mem2_26_16,
         p_wishbone_bd_ram_mem2_26_17, p_wishbone_bd_ram_mem2_26_18,
         p_wishbone_bd_ram_mem2_26_19, p_wishbone_bd_ram_mem2_26_20,
         p_wishbone_bd_ram_mem2_26_21, p_wishbone_bd_ram_mem2_26_22,
         p_wishbone_bd_ram_mem2_26_23, p_wishbone_bd_ram_mem2_27_16,
         p_wishbone_bd_ram_mem2_27_17, p_wishbone_bd_ram_mem2_27_18,
         p_wishbone_bd_ram_mem2_27_19, p_wishbone_bd_ram_mem2_27_20,
         p_wishbone_bd_ram_mem2_27_21, p_wishbone_bd_ram_mem2_27_22,
         p_wishbone_bd_ram_mem2_27_23, p_wishbone_bd_ram_mem2_28_16,
         p_wishbone_bd_ram_mem2_28_17, p_wishbone_bd_ram_mem2_28_18,
         p_wishbone_bd_ram_mem2_28_19, p_wishbone_bd_ram_mem2_28_20,
         p_wishbone_bd_ram_mem2_28_21, p_wishbone_bd_ram_mem2_28_22,
         p_wishbone_bd_ram_mem2_28_23, p_wishbone_bd_ram_mem2_29_16,
         p_wishbone_bd_ram_mem2_29_17, p_wishbone_bd_ram_mem2_29_18,
         p_wishbone_bd_ram_mem2_29_19, p_wishbone_bd_ram_mem2_29_20,
         p_wishbone_bd_ram_mem2_29_21, p_wishbone_bd_ram_mem2_29_22,
         p_wishbone_bd_ram_mem2_29_23, p_wishbone_bd_ram_mem2_30_16,
         p_wishbone_bd_ram_mem2_30_17, p_wishbone_bd_ram_mem2_30_18,
         p_wishbone_bd_ram_mem2_30_19, p_wishbone_bd_ram_mem2_30_20,
         p_wishbone_bd_ram_mem2_30_21, p_wishbone_bd_ram_mem2_30_22,
         p_wishbone_bd_ram_mem2_30_23, p_wishbone_bd_ram_mem2_31_16,
         p_wishbone_bd_ram_mem2_31_17, p_wishbone_bd_ram_mem2_31_18,
         p_wishbone_bd_ram_mem2_31_19, p_wishbone_bd_ram_mem2_31_20,
         p_wishbone_bd_ram_mem2_31_21, p_wishbone_bd_ram_mem2_31_22,
         p_wishbone_bd_ram_mem2_31_23, p_wishbone_bd_ram_mem2_32_16,
         p_wishbone_bd_ram_mem2_32_17, p_wishbone_bd_ram_mem2_32_18,
         p_wishbone_bd_ram_mem2_32_19, p_wishbone_bd_ram_mem2_32_20,
         p_wishbone_bd_ram_mem2_32_21, p_wishbone_bd_ram_mem2_32_22,
         p_wishbone_bd_ram_mem2_32_23, p_wishbone_bd_ram_mem2_33_16,
         p_wishbone_bd_ram_mem2_33_17, p_wishbone_bd_ram_mem2_33_18,
         p_wishbone_bd_ram_mem2_33_19, p_wishbone_bd_ram_mem2_33_20,
         p_wishbone_bd_ram_mem2_33_21, p_wishbone_bd_ram_mem2_33_22,
         p_wishbone_bd_ram_mem2_33_23, p_wishbone_bd_ram_mem2_34_16,
         p_wishbone_bd_ram_mem2_34_17, p_wishbone_bd_ram_mem2_34_18,
         p_wishbone_bd_ram_mem2_34_19, p_wishbone_bd_ram_mem2_34_20,
         p_wishbone_bd_ram_mem2_34_21, p_wishbone_bd_ram_mem2_34_22,
         p_wishbone_bd_ram_mem2_34_23, p_wishbone_bd_ram_mem2_35_16,
         p_wishbone_bd_ram_mem2_35_17, p_wishbone_bd_ram_mem2_35_18,
         p_wishbone_bd_ram_mem2_35_19, p_wishbone_bd_ram_mem2_35_20,
         p_wishbone_bd_ram_mem2_35_21, p_wishbone_bd_ram_mem2_35_22,
         p_wishbone_bd_ram_mem2_35_23, p_wishbone_bd_ram_mem2_36_16,
         p_wishbone_bd_ram_mem2_36_17, p_wishbone_bd_ram_mem2_36_18,
         p_wishbone_bd_ram_mem2_36_19, p_wishbone_bd_ram_mem2_36_20,
         p_wishbone_bd_ram_mem2_36_21, p_wishbone_bd_ram_mem2_36_22,
         p_wishbone_bd_ram_mem2_36_23, p_wishbone_bd_ram_mem2_37_16,
         p_wishbone_bd_ram_mem2_37_17, p_wishbone_bd_ram_mem2_37_18,
         p_wishbone_bd_ram_mem2_37_19, p_wishbone_bd_ram_mem2_37_20,
         p_wishbone_bd_ram_mem2_37_21, p_wishbone_bd_ram_mem2_37_22,
         p_wishbone_bd_ram_mem2_37_23, p_wishbone_bd_ram_mem2_38_16,
         p_wishbone_bd_ram_mem2_38_17, p_wishbone_bd_ram_mem2_38_18,
         p_wishbone_bd_ram_mem2_38_19, p_wishbone_bd_ram_mem2_38_20,
         p_wishbone_bd_ram_mem2_38_21, p_wishbone_bd_ram_mem2_38_22,
         p_wishbone_bd_ram_mem2_38_23, p_wishbone_bd_ram_mem2_39_16,
         p_wishbone_bd_ram_mem2_39_17, p_wishbone_bd_ram_mem2_39_18,
         p_wishbone_bd_ram_mem2_39_19, p_wishbone_bd_ram_mem2_39_20,
         p_wishbone_bd_ram_mem2_39_21, p_wishbone_bd_ram_mem2_39_22,
         p_wishbone_bd_ram_mem2_39_23, p_wishbone_bd_ram_mem2_40_16,
         p_wishbone_bd_ram_mem2_40_17, p_wishbone_bd_ram_mem2_40_18,
         p_wishbone_bd_ram_mem2_40_19, p_wishbone_bd_ram_mem2_40_20,
         p_wishbone_bd_ram_mem2_40_21, p_wishbone_bd_ram_mem2_40_22,
         p_wishbone_bd_ram_mem2_40_23, p_wishbone_bd_ram_mem2_41_16,
         p_wishbone_bd_ram_mem2_41_17, p_wishbone_bd_ram_mem2_41_18,
         p_wishbone_bd_ram_mem2_41_19, p_wishbone_bd_ram_mem2_41_20,
         p_wishbone_bd_ram_mem2_41_21, p_wishbone_bd_ram_mem2_41_22,
         p_wishbone_bd_ram_mem2_41_23, p_wishbone_bd_ram_mem2_42_16,
         p_wishbone_bd_ram_mem2_42_17, p_wishbone_bd_ram_mem2_42_18,
         p_wishbone_bd_ram_mem2_42_19, p_wishbone_bd_ram_mem2_42_20,
         p_wishbone_bd_ram_mem2_42_21, p_wishbone_bd_ram_mem2_42_22,
         p_wishbone_bd_ram_mem2_42_23, p_wishbone_bd_ram_mem2_43_16,
         p_wishbone_bd_ram_mem2_43_17, p_wishbone_bd_ram_mem2_43_18,
         p_wishbone_bd_ram_mem2_43_19, p_wishbone_bd_ram_mem2_43_20,
         p_wishbone_bd_ram_mem2_43_21, p_wishbone_bd_ram_mem2_43_22,
         p_wishbone_bd_ram_mem2_43_23, p_wishbone_bd_ram_mem2_44_16,
         p_wishbone_bd_ram_mem2_44_17, p_wishbone_bd_ram_mem2_44_18,
         p_wishbone_bd_ram_mem2_44_19, p_wishbone_bd_ram_mem2_44_20,
         p_wishbone_bd_ram_mem2_44_21, p_wishbone_bd_ram_mem2_44_22,
         p_wishbone_bd_ram_mem2_44_23, p_wishbone_bd_ram_mem2_45_16,
         p_wishbone_bd_ram_mem2_45_17, p_wishbone_bd_ram_mem2_45_18,
         p_wishbone_bd_ram_mem2_45_19, p_wishbone_bd_ram_mem2_45_20,
         p_wishbone_bd_ram_mem2_45_21, p_wishbone_bd_ram_mem2_45_22,
         p_wishbone_bd_ram_mem2_45_23, p_wishbone_bd_ram_mem2_46_16,
         p_wishbone_bd_ram_mem2_46_17, p_wishbone_bd_ram_mem2_46_18,
         p_wishbone_bd_ram_mem2_46_19, p_wishbone_bd_ram_mem2_46_20,
         p_wishbone_bd_ram_mem2_46_21, p_wishbone_bd_ram_mem2_46_22,
         p_wishbone_bd_ram_mem2_46_23, p_wishbone_bd_ram_mem2_47_16,
         p_wishbone_bd_ram_mem2_47_17, p_wishbone_bd_ram_mem2_47_18,
         p_wishbone_bd_ram_mem2_47_19, p_wishbone_bd_ram_mem2_47_20,
         p_wishbone_bd_ram_mem2_47_21, p_wishbone_bd_ram_mem2_47_22,
         p_wishbone_bd_ram_mem2_47_23, p_wishbone_bd_ram_mem2_48_16,
         p_wishbone_bd_ram_mem2_48_17, p_wishbone_bd_ram_mem2_48_18,
         p_wishbone_bd_ram_mem2_48_19, p_wishbone_bd_ram_mem2_48_20,
         p_wishbone_bd_ram_mem2_48_21, p_wishbone_bd_ram_mem2_48_22,
         p_wishbone_bd_ram_mem2_48_23, p_wishbone_bd_ram_mem2_49_16,
         p_wishbone_bd_ram_mem2_49_17, p_wishbone_bd_ram_mem2_49_18,
         p_wishbone_bd_ram_mem2_49_19, p_wishbone_bd_ram_mem2_49_20,
         p_wishbone_bd_ram_mem2_49_21, p_wishbone_bd_ram_mem2_49_22,
         p_wishbone_bd_ram_mem2_49_23, p_wishbone_bd_ram_mem2_50_16,
         p_wishbone_bd_ram_mem2_50_17, p_wishbone_bd_ram_mem2_50_18,
         p_wishbone_bd_ram_mem2_50_19, p_wishbone_bd_ram_mem2_50_20,
         p_wishbone_bd_ram_mem2_50_21, p_wishbone_bd_ram_mem2_50_22,
         p_wishbone_bd_ram_mem2_50_23, p_wishbone_bd_ram_mem2_51_16,
         p_wishbone_bd_ram_mem2_51_17, p_wishbone_bd_ram_mem2_51_18,
         p_wishbone_bd_ram_mem2_51_19, p_wishbone_bd_ram_mem2_51_20,
         p_wishbone_bd_ram_mem2_51_21, p_wishbone_bd_ram_mem2_51_22,
         p_wishbone_bd_ram_mem2_51_23, p_wishbone_bd_ram_mem2_52_16,
         p_wishbone_bd_ram_mem2_52_17, p_wishbone_bd_ram_mem2_52_18,
         p_wishbone_bd_ram_mem2_52_19, p_wishbone_bd_ram_mem2_52_20,
         p_wishbone_bd_ram_mem2_52_21, p_wishbone_bd_ram_mem2_52_22,
         p_wishbone_bd_ram_mem2_52_23, p_wishbone_bd_ram_mem2_53_16,
         p_wishbone_bd_ram_mem2_53_17, p_wishbone_bd_ram_mem2_53_18,
         p_wishbone_bd_ram_mem2_53_19, p_wishbone_bd_ram_mem2_53_20,
         p_wishbone_bd_ram_mem2_53_21, p_wishbone_bd_ram_mem2_53_22,
         p_wishbone_bd_ram_mem2_53_23, p_wishbone_bd_ram_mem2_54_16,
         p_wishbone_bd_ram_mem2_54_17, p_wishbone_bd_ram_mem2_54_18,
         p_wishbone_bd_ram_mem2_54_19, p_wishbone_bd_ram_mem2_54_20,
         p_wishbone_bd_ram_mem2_54_21, p_wishbone_bd_ram_mem2_54_22,
         p_wishbone_bd_ram_mem2_54_23, p_wishbone_bd_ram_mem2_55_16,
         p_wishbone_bd_ram_mem2_55_17, p_wishbone_bd_ram_mem2_55_18,
         p_wishbone_bd_ram_mem2_55_19, p_wishbone_bd_ram_mem2_55_20,
         p_wishbone_bd_ram_mem2_55_21, p_wishbone_bd_ram_mem2_55_22,
         p_wishbone_bd_ram_mem2_55_23, p_wishbone_bd_ram_mem2_56_16,
         p_wishbone_bd_ram_mem2_56_17, p_wishbone_bd_ram_mem2_56_18,
         p_wishbone_bd_ram_mem2_56_19, p_wishbone_bd_ram_mem2_56_20,
         p_wishbone_bd_ram_mem2_56_21, p_wishbone_bd_ram_mem2_56_22,
         p_wishbone_bd_ram_mem2_56_23, p_wishbone_bd_ram_mem2_57_16,
         p_wishbone_bd_ram_mem2_57_17, p_wishbone_bd_ram_mem2_57_18,
         p_wishbone_bd_ram_mem2_57_19, p_wishbone_bd_ram_mem2_57_20,
         p_wishbone_bd_ram_mem2_57_21, p_wishbone_bd_ram_mem2_57_22,
         p_wishbone_bd_ram_mem2_57_23, p_wishbone_bd_ram_mem2_58_16,
         p_wishbone_bd_ram_mem2_58_17, p_wishbone_bd_ram_mem2_58_18,
         p_wishbone_bd_ram_mem2_58_19, p_wishbone_bd_ram_mem2_58_20,
         p_wishbone_bd_ram_mem2_58_21, p_wishbone_bd_ram_mem2_58_22,
         p_wishbone_bd_ram_mem2_58_23, p_wishbone_bd_ram_mem2_59_16,
         p_wishbone_bd_ram_mem2_59_17, p_wishbone_bd_ram_mem2_59_18,
         p_wishbone_bd_ram_mem2_59_19, p_wishbone_bd_ram_mem2_59_20,
         p_wishbone_bd_ram_mem2_59_21, p_wishbone_bd_ram_mem2_59_22,
         p_wishbone_bd_ram_mem2_59_23, p_wishbone_bd_ram_mem2_60_16,
         p_wishbone_bd_ram_mem2_60_17, p_wishbone_bd_ram_mem2_60_18,
         p_wishbone_bd_ram_mem2_60_19, p_wishbone_bd_ram_mem2_60_20,
         p_wishbone_bd_ram_mem2_60_21, p_wishbone_bd_ram_mem2_60_22,
         p_wishbone_bd_ram_mem2_60_23, p_wishbone_bd_ram_mem2_61_16,
         p_wishbone_bd_ram_mem2_61_17, p_wishbone_bd_ram_mem2_61_18,
         p_wishbone_bd_ram_mem2_61_19, p_wishbone_bd_ram_mem2_61_20,
         p_wishbone_bd_ram_mem2_61_21, p_wishbone_bd_ram_mem2_61_22,
         p_wishbone_bd_ram_mem2_61_23, p_wishbone_bd_ram_mem2_62_16,
         p_wishbone_bd_ram_mem2_62_17, p_wishbone_bd_ram_mem2_62_18,
         p_wishbone_bd_ram_mem2_62_19, p_wishbone_bd_ram_mem2_62_20,
         p_wishbone_bd_ram_mem2_62_21, p_wishbone_bd_ram_mem2_62_22,
         p_wishbone_bd_ram_mem2_62_23, p_wishbone_bd_ram_mem2_63_16,
         p_wishbone_bd_ram_mem2_63_17, p_wishbone_bd_ram_mem2_63_18,
         p_wishbone_bd_ram_mem2_63_19, p_wishbone_bd_ram_mem2_63_20,
         p_wishbone_bd_ram_mem2_63_21, p_wishbone_bd_ram_mem2_63_22,
         p_wishbone_bd_ram_mem2_63_23, p_wishbone_bd_ram_mem2_64_16,
         p_wishbone_bd_ram_mem2_64_17, p_wishbone_bd_ram_mem2_64_18,
         p_wishbone_bd_ram_mem2_64_19, p_wishbone_bd_ram_mem2_64_20,
         p_wishbone_bd_ram_mem2_64_21, p_wishbone_bd_ram_mem2_64_22,
         p_wishbone_bd_ram_mem2_64_23, p_wishbone_bd_ram_mem2_65_16,
         p_wishbone_bd_ram_mem2_65_17, p_wishbone_bd_ram_mem2_65_18,
         p_wishbone_bd_ram_mem2_65_19, p_wishbone_bd_ram_mem2_65_20,
         p_wishbone_bd_ram_mem2_65_21, p_wishbone_bd_ram_mem2_65_22,
         p_wishbone_bd_ram_mem2_65_23, p_wishbone_bd_ram_mem2_66_16,
         p_wishbone_bd_ram_mem2_66_17, p_wishbone_bd_ram_mem2_66_18,
         p_wishbone_bd_ram_mem2_66_19, p_wishbone_bd_ram_mem2_66_20,
         p_wishbone_bd_ram_mem2_66_21, p_wishbone_bd_ram_mem2_66_22,
         p_wishbone_bd_ram_mem2_66_23, p_wishbone_bd_ram_mem2_67_16,
         p_wishbone_bd_ram_mem2_67_17, p_wishbone_bd_ram_mem2_67_18,
         p_wishbone_bd_ram_mem2_67_19, p_wishbone_bd_ram_mem2_67_20,
         p_wishbone_bd_ram_mem2_67_21, p_wishbone_bd_ram_mem2_67_22,
         p_wishbone_bd_ram_mem2_67_23, p_wishbone_bd_ram_mem2_68_16,
         p_wishbone_bd_ram_mem2_68_17, p_wishbone_bd_ram_mem2_68_18,
         p_wishbone_bd_ram_mem2_68_19, p_wishbone_bd_ram_mem2_68_20,
         p_wishbone_bd_ram_mem2_68_21, p_wishbone_bd_ram_mem2_68_22,
         p_wishbone_bd_ram_mem2_68_23, p_wishbone_bd_ram_mem2_69_16,
         p_wishbone_bd_ram_mem2_69_17, p_wishbone_bd_ram_mem2_69_18,
         p_wishbone_bd_ram_mem2_69_19, p_wishbone_bd_ram_mem2_69_20,
         p_wishbone_bd_ram_mem2_69_21, p_wishbone_bd_ram_mem2_69_22,
         p_wishbone_bd_ram_mem2_69_23, p_wishbone_bd_ram_mem2_70_16,
         p_wishbone_bd_ram_mem2_70_17, p_wishbone_bd_ram_mem2_70_18,
         p_wishbone_bd_ram_mem2_70_19, p_wishbone_bd_ram_mem2_70_20,
         p_wishbone_bd_ram_mem2_70_21, p_wishbone_bd_ram_mem2_70_22,
         p_wishbone_bd_ram_mem2_70_23, p_wishbone_bd_ram_mem2_71_16,
         p_wishbone_bd_ram_mem2_71_17, p_wishbone_bd_ram_mem2_71_18,
         p_wishbone_bd_ram_mem2_71_19, p_wishbone_bd_ram_mem2_71_20,
         p_wishbone_bd_ram_mem2_71_21, p_wishbone_bd_ram_mem2_71_22,
         p_wishbone_bd_ram_mem2_71_23, p_wishbone_bd_ram_mem2_72_16,
         p_wishbone_bd_ram_mem2_72_17, p_wishbone_bd_ram_mem2_72_18,
         p_wishbone_bd_ram_mem2_72_19, p_wishbone_bd_ram_mem2_72_20,
         p_wishbone_bd_ram_mem2_72_21, p_wishbone_bd_ram_mem2_72_22,
         p_wishbone_bd_ram_mem2_72_23, p_wishbone_bd_ram_mem2_73_16,
         p_wishbone_bd_ram_mem2_73_17, p_wishbone_bd_ram_mem2_73_18,
         p_wishbone_bd_ram_mem2_73_19, p_wishbone_bd_ram_mem2_73_20,
         p_wishbone_bd_ram_mem2_73_21, p_wishbone_bd_ram_mem2_73_22,
         p_wishbone_bd_ram_mem2_73_23, p_wishbone_bd_ram_mem2_74_16,
         p_wishbone_bd_ram_mem2_74_17, p_wishbone_bd_ram_mem2_74_18,
         p_wishbone_bd_ram_mem2_74_19, p_wishbone_bd_ram_mem2_74_20,
         p_wishbone_bd_ram_mem2_74_21, p_wishbone_bd_ram_mem2_74_22,
         p_wishbone_bd_ram_mem2_74_23, p_wishbone_bd_ram_mem2_75_16,
         p_wishbone_bd_ram_mem2_75_17, p_wishbone_bd_ram_mem2_75_18,
         p_wishbone_bd_ram_mem2_75_19, p_wishbone_bd_ram_mem2_75_20,
         p_wishbone_bd_ram_mem2_75_21, p_wishbone_bd_ram_mem2_75_22,
         p_wishbone_bd_ram_mem2_75_23, p_wishbone_bd_ram_mem2_76_16,
         p_wishbone_bd_ram_mem2_76_17, p_wishbone_bd_ram_mem2_76_18,
         p_wishbone_bd_ram_mem2_76_19, p_wishbone_bd_ram_mem2_76_20,
         p_wishbone_bd_ram_mem2_76_21, p_wishbone_bd_ram_mem2_76_22,
         p_wishbone_bd_ram_mem2_76_23, p_wishbone_bd_ram_mem2_77_16,
         p_wishbone_bd_ram_mem2_77_17, p_wishbone_bd_ram_mem2_77_18,
         p_wishbone_bd_ram_mem2_77_19, p_wishbone_bd_ram_mem2_77_20,
         p_wishbone_bd_ram_mem2_77_21, p_wishbone_bd_ram_mem2_77_22,
         p_wishbone_bd_ram_mem2_77_23, p_wishbone_bd_ram_mem2_78_16,
         p_wishbone_bd_ram_mem2_78_17, p_wishbone_bd_ram_mem2_78_18,
         p_wishbone_bd_ram_mem2_78_19, p_wishbone_bd_ram_mem2_78_20,
         p_wishbone_bd_ram_mem2_78_21, p_wishbone_bd_ram_mem2_78_22,
         p_wishbone_bd_ram_mem2_78_23, p_wishbone_bd_ram_mem2_79_16,
         p_wishbone_bd_ram_mem2_79_17, p_wishbone_bd_ram_mem2_79_18,
         p_wishbone_bd_ram_mem2_79_19, p_wishbone_bd_ram_mem2_79_20,
         p_wishbone_bd_ram_mem2_79_21, p_wishbone_bd_ram_mem2_79_22,
         p_wishbone_bd_ram_mem2_79_23, p_wishbone_bd_ram_mem2_80_16,
         p_wishbone_bd_ram_mem2_80_17, p_wishbone_bd_ram_mem2_80_18,
         p_wishbone_bd_ram_mem2_80_19, p_wishbone_bd_ram_mem2_80_20,
         p_wishbone_bd_ram_mem2_80_21, p_wishbone_bd_ram_mem2_80_22,
         p_wishbone_bd_ram_mem2_80_23, p_wishbone_bd_ram_mem2_81_16,
         p_wishbone_bd_ram_mem2_81_17, p_wishbone_bd_ram_mem2_81_18,
         p_wishbone_bd_ram_mem2_81_19, p_wishbone_bd_ram_mem2_81_20,
         p_wishbone_bd_ram_mem2_81_21, p_wishbone_bd_ram_mem2_81_22,
         p_wishbone_bd_ram_mem2_81_23, p_wishbone_bd_ram_mem2_82_16,
         p_wishbone_bd_ram_mem2_82_17, p_wishbone_bd_ram_mem2_82_18,
         p_wishbone_bd_ram_mem2_82_19, p_wishbone_bd_ram_mem2_82_20,
         p_wishbone_bd_ram_mem2_82_21, p_wishbone_bd_ram_mem2_82_22,
         p_wishbone_bd_ram_mem2_82_23, p_wishbone_bd_ram_mem2_83_16,
         p_wishbone_bd_ram_mem2_83_17, p_wishbone_bd_ram_mem2_83_18,
         p_wishbone_bd_ram_mem2_83_19, p_wishbone_bd_ram_mem2_83_20,
         p_wishbone_bd_ram_mem2_83_21, p_wishbone_bd_ram_mem2_83_22,
         p_wishbone_bd_ram_mem2_83_23, p_wishbone_bd_ram_mem2_84_16,
         p_wishbone_bd_ram_mem2_84_17, p_wishbone_bd_ram_mem2_84_18,
         p_wishbone_bd_ram_mem2_84_19, p_wishbone_bd_ram_mem2_84_20,
         p_wishbone_bd_ram_mem2_84_21, p_wishbone_bd_ram_mem2_84_22,
         p_wishbone_bd_ram_mem2_84_23, p_wishbone_bd_ram_mem2_85_16,
         p_wishbone_bd_ram_mem2_85_17, p_wishbone_bd_ram_mem2_85_18,
         p_wishbone_bd_ram_mem2_85_19, p_wishbone_bd_ram_mem2_85_20,
         p_wishbone_bd_ram_mem2_85_21, p_wishbone_bd_ram_mem2_85_22,
         p_wishbone_bd_ram_mem2_85_23, p_wishbone_bd_ram_mem2_86_16,
         p_wishbone_bd_ram_mem2_86_17, p_wishbone_bd_ram_mem2_86_18,
         p_wishbone_bd_ram_mem2_86_19, p_wishbone_bd_ram_mem2_86_20,
         p_wishbone_bd_ram_mem2_86_21, p_wishbone_bd_ram_mem2_86_22,
         p_wishbone_bd_ram_mem2_86_23, p_wishbone_bd_ram_mem2_87_16,
         p_wishbone_bd_ram_mem2_87_17, p_wishbone_bd_ram_mem2_87_18,
         p_wishbone_bd_ram_mem2_87_19, p_wishbone_bd_ram_mem2_87_20,
         p_wishbone_bd_ram_mem2_87_21, p_wishbone_bd_ram_mem2_87_22,
         p_wishbone_bd_ram_mem2_87_23, p_wishbone_bd_ram_mem2_88_16,
         p_wishbone_bd_ram_mem2_88_17, p_wishbone_bd_ram_mem2_88_18,
         p_wishbone_bd_ram_mem2_88_19, p_wishbone_bd_ram_mem2_88_20,
         p_wishbone_bd_ram_mem2_88_21, p_wishbone_bd_ram_mem2_88_22,
         p_wishbone_bd_ram_mem2_88_23, p_wishbone_bd_ram_mem2_89_16,
         p_wishbone_bd_ram_mem2_89_17, p_wishbone_bd_ram_mem2_89_18,
         p_wishbone_bd_ram_mem2_89_19, p_wishbone_bd_ram_mem2_89_20,
         p_wishbone_bd_ram_mem2_89_21, p_wishbone_bd_ram_mem2_89_22,
         p_wishbone_bd_ram_mem2_89_23, p_wishbone_bd_ram_mem2_90_16,
         p_wishbone_bd_ram_mem2_90_17, p_wishbone_bd_ram_mem2_90_18,
         p_wishbone_bd_ram_mem2_90_19, p_wishbone_bd_ram_mem2_90_20,
         p_wishbone_bd_ram_mem2_90_21, p_wishbone_bd_ram_mem2_90_22,
         p_wishbone_bd_ram_mem2_90_23, p_wishbone_bd_ram_mem2_91_16,
         p_wishbone_bd_ram_mem2_91_17, p_wishbone_bd_ram_mem2_91_18,
         p_wishbone_bd_ram_mem2_91_19, p_wishbone_bd_ram_mem2_91_20,
         p_wishbone_bd_ram_mem2_91_21, p_wishbone_bd_ram_mem2_91_22,
         p_wishbone_bd_ram_mem2_91_23, p_wishbone_bd_ram_mem2_92_16,
         p_wishbone_bd_ram_mem2_92_17, p_wishbone_bd_ram_mem2_92_18,
         p_wishbone_bd_ram_mem2_92_19, p_wishbone_bd_ram_mem2_92_20,
         p_wishbone_bd_ram_mem2_92_21, p_wishbone_bd_ram_mem2_92_22,
         p_wishbone_bd_ram_mem2_92_23, p_wishbone_bd_ram_mem2_93_16,
         p_wishbone_bd_ram_mem2_93_17, p_wishbone_bd_ram_mem2_93_18,
         p_wishbone_bd_ram_mem2_93_19, p_wishbone_bd_ram_mem2_93_20,
         p_wishbone_bd_ram_mem2_93_21, p_wishbone_bd_ram_mem2_93_22,
         p_wishbone_bd_ram_mem2_93_23, p_wishbone_bd_ram_mem2_94_16,
         p_wishbone_bd_ram_mem2_94_17, p_wishbone_bd_ram_mem2_94_18,
         p_wishbone_bd_ram_mem2_94_19, p_wishbone_bd_ram_mem2_94_20,
         p_wishbone_bd_ram_mem2_94_21, p_wishbone_bd_ram_mem2_94_22,
         p_wishbone_bd_ram_mem2_94_23, p_wishbone_bd_ram_mem2_95_16,
         p_wishbone_bd_ram_mem2_95_17, p_wishbone_bd_ram_mem2_95_18,
         p_wishbone_bd_ram_mem2_95_19, p_wishbone_bd_ram_mem2_95_20,
         p_wishbone_bd_ram_mem2_95_21, p_wishbone_bd_ram_mem2_95_22,
         p_wishbone_bd_ram_mem2_95_23, p_wishbone_bd_ram_mem2_96_16,
         p_wishbone_bd_ram_mem2_96_17, p_wishbone_bd_ram_mem2_96_18,
         p_wishbone_bd_ram_mem2_96_19, p_wishbone_bd_ram_mem2_96_20,
         p_wishbone_bd_ram_mem2_96_21, p_wishbone_bd_ram_mem2_96_22,
         p_wishbone_bd_ram_mem2_96_23, p_wishbone_bd_ram_mem2_97_16,
         p_wishbone_bd_ram_mem2_97_17, p_wishbone_bd_ram_mem2_97_18,
         p_wishbone_bd_ram_mem2_97_19, p_wishbone_bd_ram_mem2_97_20,
         p_wishbone_bd_ram_mem2_97_21, p_wishbone_bd_ram_mem2_97_22,
         p_wishbone_bd_ram_mem2_97_23, p_wishbone_bd_ram_mem2_98_16,
         p_wishbone_bd_ram_mem2_98_17, p_wishbone_bd_ram_mem2_98_18,
         p_wishbone_bd_ram_mem2_98_19, p_wishbone_bd_ram_mem2_98_20,
         p_wishbone_bd_ram_mem2_98_21, p_wishbone_bd_ram_mem2_98_22,
         p_wishbone_bd_ram_mem2_98_23, p_wishbone_bd_ram_mem2_99_16,
         p_wishbone_bd_ram_mem2_99_17, p_wishbone_bd_ram_mem2_99_18,
         p_wishbone_bd_ram_mem2_99_19, p_wishbone_bd_ram_mem2_99_20,
         p_wishbone_bd_ram_mem2_99_21, p_wishbone_bd_ram_mem2_99_22,
         p_wishbone_bd_ram_mem2_99_23, p_wishbone_bd_ram_mem2_100_16,
         p_wishbone_bd_ram_mem2_100_17, p_wishbone_bd_ram_mem2_100_18,
         p_wishbone_bd_ram_mem2_100_19, p_wishbone_bd_ram_mem2_100_20,
         p_wishbone_bd_ram_mem2_100_21, p_wishbone_bd_ram_mem2_100_22,
         p_wishbone_bd_ram_mem2_100_23, p_wishbone_bd_ram_mem2_101_16,
         p_wishbone_bd_ram_mem2_101_17, p_wishbone_bd_ram_mem2_101_18,
         p_wishbone_bd_ram_mem2_101_19, p_wishbone_bd_ram_mem2_101_20,
         p_wishbone_bd_ram_mem2_101_21, p_wishbone_bd_ram_mem2_101_22,
         p_wishbone_bd_ram_mem2_101_23, p_wishbone_bd_ram_mem2_102_16,
         p_wishbone_bd_ram_mem2_102_17, p_wishbone_bd_ram_mem2_102_18,
         p_wishbone_bd_ram_mem2_102_19, p_wishbone_bd_ram_mem2_102_20,
         p_wishbone_bd_ram_mem2_102_21, p_wishbone_bd_ram_mem2_102_22,
         p_wishbone_bd_ram_mem2_102_23, p_wishbone_bd_ram_mem2_103_16,
         p_wishbone_bd_ram_mem2_103_17, p_wishbone_bd_ram_mem2_103_18,
         p_wishbone_bd_ram_mem2_103_19, p_wishbone_bd_ram_mem2_103_20,
         p_wishbone_bd_ram_mem2_103_21, p_wishbone_bd_ram_mem2_103_22,
         p_wishbone_bd_ram_mem2_103_23, p_wishbone_bd_ram_mem2_104_16,
         p_wishbone_bd_ram_mem2_104_17, p_wishbone_bd_ram_mem2_104_18,
         p_wishbone_bd_ram_mem2_104_19, p_wishbone_bd_ram_mem2_104_20,
         p_wishbone_bd_ram_mem2_104_21, p_wishbone_bd_ram_mem2_104_22,
         p_wishbone_bd_ram_mem2_104_23, p_wishbone_bd_ram_mem2_105_16,
         p_wishbone_bd_ram_mem2_105_17, p_wishbone_bd_ram_mem2_105_18,
         p_wishbone_bd_ram_mem2_105_19, p_wishbone_bd_ram_mem2_105_20,
         p_wishbone_bd_ram_mem2_105_21, p_wishbone_bd_ram_mem2_105_22,
         p_wishbone_bd_ram_mem2_105_23, p_wishbone_bd_ram_mem2_106_16,
         p_wishbone_bd_ram_mem2_106_17, p_wishbone_bd_ram_mem2_106_18,
         p_wishbone_bd_ram_mem2_106_19, p_wishbone_bd_ram_mem2_106_20,
         p_wishbone_bd_ram_mem2_106_21, p_wishbone_bd_ram_mem2_106_22,
         p_wishbone_bd_ram_mem2_106_23, p_wishbone_bd_ram_mem2_107_16,
         p_wishbone_bd_ram_mem2_107_17, p_wishbone_bd_ram_mem2_107_18,
         p_wishbone_bd_ram_mem2_107_19, p_wishbone_bd_ram_mem2_107_20,
         p_wishbone_bd_ram_mem2_107_21, p_wishbone_bd_ram_mem2_107_22,
         p_wishbone_bd_ram_mem2_107_23, p_wishbone_bd_ram_mem2_108_16,
         p_wishbone_bd_ram_mem2_108_17, p_wishbone_bd_ram_mem2_108_18,
         p_wishbone_bd_ram_mem2_108_19, p_wishbone_bd_ram_mem2_108_20,
         p_wishbone_bd_ram_mem2_108_21, p_wishbone_bd_ram_mem2_108_22,
         p_wishbone_bd_ram_mem2_108_23, p_wishbone_bd_ram_mem2_109_16,
         p_wishbone_bd_ram_mem2_109_17, p_wishbone_bd_ram_mem2_109_18,
         p_wishbone_bd_ram_mem2_109_19, p_wishbone_bd_ram_mem2_109_20,
         p_wishbone_bd_ram_mem2_109_21, p_wishbone_bd_ram_mem2_109_22,
         p_wishbone_bd_ram_mem2_109_23, p_wishbone_bd_ram_mem2_110_16,
         p_wishbone_bd_ram_mem2_110_17, p_wishbone_bd_ram_mem2_110_18,
         p_wishbone_bd_ram_mem2_110_19, p_wishbone_bd_ram_mem2_110_20,
         p_wishbone_bd_ram_mem2_110_21, p_wishbone_bd_ram_mem2_110_22,
         p_wishbone_bd_ram_mem2_110_23, p_wishbone_bd_ram_mem2_111_16,
         p_wishbone_bd_ram_mem2_111_17, p_wishbone_bd_ram_mem2_111_18,
         p_wishbone_bd_ram_mem2_111_19, p_wishbone_bd_ram_mem2_111_20,
         p_wishbone_bd_ram_mem2_111_21, p_wishbone_bd_ram_mem2_111_22,
         p_wishbone_bd_ram_mem2_111_23, p_wishbone_bd_ram_mem2_112_16,
         p_wishbone_bd_ram_mem2_112_17, p_wishbone_bd_ram_mem2_112_18,
         p_wishbone_bd_ram_mem2_112_19, p_wishbone_bd_ram_mem2_112_20,
         p_wishbone_bd_ram_mem2_112_21, p_wishbone_bd_ram_mem2_112_22,
         p_wishbone_bd_ram_mem2_112_23, p_wishbone_bd_ram_mem2_113_16,
         p_wishbone_bd_ram_mem2_113_17, p_wishbone_bd_ram_mem2_113_18,
         p_wishbone_bd_ram_mem2_113_19, p_wishbone_bd_ram_mem2_113_20,
         p_wishbone_bd_ram_mem2_113_21, p_wishbone_bd_ram_mem2_113_22,
         p_wishbone_bd_ram_mem2_113_23, p_wishbone_bd_ram_mem2_114_16,
         p_wishbone_bd_ram_mem2_114_17, p_wishbone_bd_ram_mem2_114_18,
         p_wishbone_bd_ram_mem2_114_19, p_wishbone_bd_ram_mem2_114_20,
         p_wishbone_bd_ram_mem2_114_21, p_wishbone_bd_ram_mem2_114_22,
         p_wishbone_bd_ram_mem2_114_23, p_wishbone_bd_ram_mem2_115_16,
         p_wishbone_bd_ram_mem2_115_17, p_wishbone_bd_ram_mem2_115_18,
         p_wishbone_bd_ram_mem2_115_19, p_wishbone_bd_ram_mem2_115_20,
         p_wishbone_bd_ram_mem2_115_21, p_wishbone_bd_ram_mem2_115_22,
         p_wishbone_bd_ram_mem2_115_23, p_wishbone_bd_ram_mem2_116_16,
         p_wishbone_bd_ram_mem2_116_17, p_wishbone_bd_ram_mem2_116_18,
         p_wishbone_bd_ram_mem2_116_19, p_wishbone_bd_ram_mem2_116_20,
         p_wishbone_bd_ram_mem2_116_21, p_wishbone_bd_ram_mem2_116_22,
         p_wishbone_bd_ram_mem2_116_23, p_wishbone_bd_ram_mem2_117_16,
         p_wishbone_bd_ram_mem2_117_17, p_wishbone_bd_ram_mem2_117_18,
         p_wishbone_bd_ram_mem2_117_19, p_wishbone_bd_ram_mem2_117_20,
         p_wishbone_bd_ram_mem2_117_21, p_wishbone_bd_ram_mem2_117_22,
         p_wishbone_bd_ram_mem2_117_23, p_wishbone_bd_ram_mem2_118_16,
         p_wishbone_bd_ram_mem2_118_17, p_wishbone_bd_ram_mem2_118_18,
         p_wishbone_bd_ram_mem2_118_19, p_wishbone_bd_ram_mem2_118_20,
         p_wishbone_bd_ram_mem2_118_21, p_wishbone_bd_ram_mem2_118_22,
         p_wishbone_bd_ram_mem2_118_23, p_wishbone_bd_ram_mem2_119_16,
         p_wishbone_bd_ram_mem2_119_17, p_wishbone_bd_ram_mem2_119_18,
         p_wishbone_bd_ram_mem2_119_19, p_wishbone_bd_ram_mem2_119_20,
         p_wishbone_bd_ram_mem2_119_21, p_wishbone_bd_ram_mem2_119_22,
         p_wishbone_bd_ram_mem2_119_23, p_wishbone_bd_ram_mem2_120_16,
         p_wishbone_bd_ram_mem2_120_17, p_wishbone_bd_ram_mem2_120_18,
         p_wishbone_bd_ram_mem2_120_19, p_wishbone_bd_ram_mem2_120_20,
         p_wishbone_bd_ram_mem2_120_21, p_wishbone_bd_ram_mem2_120_22,
         p_wishbone_bd_ram_mem2_120_23, p_wishbone_bd_ram_mem2_121_16,
         p_wishbone_bd_ram_mem2_121_17, p_wishbone_bd_ram_mem2_121_18,
         p_wishbone_bd_ram_mem2_121_19, p_wishbone_bd_ram_mem2_121_20,
         p_wishbone_bd_ram_mem2_121_21, p_wishbone_bd_ram_mem2_121_22,
         p_wishbone_bd_ram_mem2_121_23, p_wishbone_bd_ram_mem2_122_16,
         p_wishbone_bd_ram_mem2_122_17, p_wishbone_bd_ram_mem2_122_18,
         p_wishbone_bd_ram_mem2_122_19, p_wishbone_bd_ram_mem2_122_20,
         p_wishbone_bd_ram_mem2_122_21, p_wishbone_bd_ram_mem2_122_22,
         p_wishbone_bd_ram_mem2_122_23, p_wishbone_bd_ram_mem2_123_16,
         p_wishbone_bd_ram_mem2_123_17, p_wishbone_bd_ram_mem2_123_18,
         p_wishbone_bd_ram_mem2_123_19, p_wishbone_bd_ram_mem2_123_20,
         p_wishbone_bd_ram_mem2_123_21, p_wishbone_bd_ram_mem2_123_22,
         p_wishbone_bd_ram_mem2_123_23, p_wishbone_bd_ram_mem2_124_16,
         p_wishbone_bd_ram_mem2_124_17, p_wishbone_bd_ram_mem2_124_18,
         p_wishbone_bd_ram_mem2_124_19, p_wishbone_bd_ram_mem2_124_20,
         p_wishbone_bd_ram_mem2_124_21, p_wishbone_bd_ram_mem2_124_22,
         p_wishbone_bd_ram_mem2_124_23, p_wishbone_bd_ram_mem2_125_16,
         p_wishbone_bd_ram_mem2_125_17, p_wishbone_bd_ram_mem2_125_18,
         p_wishbone_bd_ram_mem2_125_19, p_wishbone_bd_ram_mem2_125_20,
         p_wishbone_bd_ram_mem2_125_21, p_wishbone_bd_ram_mem2_125_22,
         p_wishbone_bd_ram_mem2_125_23, p_wishbone_bd_ram_mem2_126_16,
         p_wishbone_bd_ram_mem2_126_17, p_wishbone_bd_ram_mem2_126_18,
         p_wishbone_bd_ram_mem2_126_19, p_wishbone_bd_ram_mem2_126_20,
         p_wishbone_bd_ram_mem2_126_21, p_wishbone_bd_ram_mem2_126_22,
         p_wishbone_bd_ram_mem2_126_23, p_wishbone_bd_ram_mem2_127_16,
         p_wishbone_bd_ram_mem2_127_17, p_wishbone_bd_ram_mem2_127_18,
         p_wishbone_bd_ram_mem2_127_19, p_wishbone_bd_ram_mem2_127_20,
         p_wishbone_bd_ram_mem2_127_21, p_wishbone_bd_ram_mem2_127_22,
         p_wishbone_bd_ram_mem2_127_23, p_wishbone_bd_ram_mem2_128_16,
         p_wishbone_bd_ram_mem2_128_17, p_wishbone_bd_ram_mem2_128_18,
         p_wishbone_bd_ram_mem2_128_19, p_wishbone_bd_ram_mem2_128_20,
         p_wishbone_bd_ram_mem2_128_21, p_wishbone_bd_ram_mem2_128_22,
         p_wishbone_bd_ram_mem2_128_23, p_wishbone_bd_ram_mem2_129_16,
         p_wishbone_bd_ram_mem2_129_17, p_wishbone_bd_ram_mem2_129_18,
         p_wishbone_bd_ram_mem2_129_19, p_wishbone_bd_ram_mem2_129_20,
         p_wishbone_bd_ram_mem2_129_21, p_wishbone_bd_ram_mem2_129_22,
         p_wishbone_bd_ram_mem2_129_23, p_wishbone_bd_ram_mem2_130_16,
         p_wishbone_bd_ram_mem2_130_17, p_wishbone_bd_ram_mem2_130_18,
         p_wishbone_bd_ram_mem2_130_19, p_wishbone_bd_ram_mem2_130_20,
         p_wishbone_bd_ram_mem2_130_21, p_wishbone_bd_ram_mem2_130_22,
         p_wishbone_bd_ram_mem2_130_23, p_wishbone_bd_ram_mem2_131_16,
         p_wishbone_bd_ram_mem2_131_17, p_wishbone_bd_ram_mem2_131_18,
         p_wishbone_bd_ram_mem2_131_19, p_wishbone_bd_ram_mem2_131_20,
         p_wishbone_bd_ram_mem2_131_21, p_wishbone_bd_ram_mem2_131_22,
         p_wishbone_bd_ram_mem2_131_23, p_wishbone_bd_ram_mem2_132_16,
         p_wishbone_bd_ram_mem2_132_17, p_wishbone_bd_ram_mem2_132_18,
         p_wishbone_bd_ram_mem2_132_19, p_wishbone_bd_ram_mem2_132_20,
         p_wishbone_bd_ram_mem2_132_21, p_wishbone_bd_ram_mem2_132_22,
         p_wishbone_bd_ram_mem2_132_23, p_wishbone_bd_ram_mem2_133_16,
         p_wishbone_bd_ram_mem2_133_17, p_wishbone_bd_ram_mem2_133_18,
         p_wishbone_bd_ram_mem2_133_19, p_wishbone_bd_ram_mem2_133_20,
         p_wishbone_bd_ram_mem2_133_21, p_wishbone_bd_ram_mem2_133_22,
         p_wishbone_bd_ram_mem2_133_23, p_wishbone_bd_ram_mem2_134_16,
         p_wishbone_bd_ram_mem2_134_17, p_wishbone_bd_ram_mem2_134_18,
         p_wishbone_bd_ram_mem2_134_19, p_wishbone_bd_ram_mem2_134_20,
         p_wishbone_bd_ram_mem2_134_21, p_wishbone_bd_ram_mem2_134_22,
         p_wishbone_bd_ram_mem2_134_23, p_wishbone_bd_ram_mem2_135_16,
         p_wishbone_bd_ram_mem2_135_17, p_wishbone_bd_ram_mem2_135_18,
         p_wishbone_bd_ram_mem2_135_19, p_wishbone_bd_ram_mem2_135_20,
         p_wishbone_bd_ram_mem2_135_21, p_wishbone_bd_ram_mem2_135_22,
         p_wishbone_bd_ram_mem2_135_23, p_wishbone_bd_ram_mem2_136_16,
         p_wishbone_bd_ram_mem2_136_17, p_wishbone_bd_ram_mem2_136_18,
         p_wishbone_bd_ram_mem2_136_19, p_wishbone_bd_ram_mem2_136_20,
         p_wishbone_bd_ram_mem2_136_21, p_wishbone_bd_ram_mem2_136_22,
         p_wishbone_bd_ram_mem2_136_23, p_wishbone_bd_ram_mem2_137_16,
         p_wishbone_bd_ram_mem2_137_17, p_wishbone_bd_ram_mem2_137_18,
         p_wishbone_bd_ram_mem2_137_19, p_wishbone_bd_ram_mem2_137_20,
         p_wishbone_bd_ram_mem2_137_21, p_wishbone_bd_ram_mem2_137_22,
         p_wishbone_bd_ram_mem2_137_23, p_wishbone_bd_ram_mem2_138_16,
         p_wishbone_bd_ram_mem2_138_17, p_wishbone_bd_ram_mem2_138_18,
         p_wishbone_bd_ram_mem2_138_19, p_wishbone_bd_ram_mem2_138_20,
         p_wishbone_bd_ram_mem2_138_21, p_wishbone_bd_ram_mem2_138_22,
         p_wishbone_bd_ram_mem2_138_23, p_wishbone_bd_ram_mem2_139_16,
         p_wishbone_bd_ram_mem2_139_17, p_wishbone_bd_ram_mem2_139_18,
         p_wishbone_bd_ram_mem2_139_19, p_wishbone_bd_ram_mem2_139_20,
         p_wishbone_bd_ram_mem2_139_21, p_wishbone_bd_ram_mem2_139_22,
         p_wishbone_bd_ram_mem2_139_23, p_wishbone_bd_ram_mem2_140_16,
         p_wishbone_bd_ram_mem2_140_17, p_wishbone_bd_ram_mem2_140_18,
         p_wishbone_bd_ram_mem2_140_19, p_wishbone_bd_ram_mem2_140_20,
         p_wishbone_bd_ram_mem2_140_21, p_wishbone_bd_ram_mem2_140_22,
         p_wishbone_bd_ram_mem2_140_23, p_wishbone_bd_ram_mem2_141_16,
         p_wishbone_bd_ram_mem2_141_17, p_wishbone_bd_ram_mem2_141_18,
         p_wishbone_bd_ram_mem2_141_19, p_wishbone_bd_ram_mem2_141_20,
         p_wishbone_bd_ram_mem2_141_21, p_wishbone_bd_ram_mem2_141_22,
         p_wishbone_bd_ram_mem2_141_23, p_wishbone_bd_ram_mem2_142_16,
         p_wishbone_bd_ram_mem2_142_17, p_wishbone_bd_ram_mem2_142_18,
         p_wishbone_bd_ram_mem2_142_19, p_wishbone_bd_ram_mem2_142_20,
         p_wishbone_bd_ram_mem2_142_21, p_wishbone_bd_ram_mem2_142_22,
         p_wishbone_bd_ram_mem2_142_23, p_wishbone_bd_ram_mem2_143_16,
         p_wishbone_bd_ram_mem2_143_17, p_wishbone_bd_ram_mem2_143_18,
         p_wishbone_bd_ram_mem2_143_19, p_wishbone_bd_ram_mem2_143_20,
         p_wishbone_bd_ram_mem2_143_21, p_wishbone_bd_ram_mem2_143_22,
         p_wishbone_bd_ram_mem2_143_23, p_wishbone_bd_ram_mem2_144_16,
         p_wishbone_bd_ram_mem2_144_17, p_wishbone_bd_ram_mem2_144_18,
         p_wishbone_bd_ram_mem2_144_19, p_wishbone_bd_ram_mem2_144_20,
         p_wishbone_bd_ram_mem2_144_21, p_wishbone_bd_ram_mem2_144_22,
         p_wishbone_bd_ram_mem2_144_23, p_wishbone_bd_ram_mem2_145_16,
         p_wishbone_bd_ram_mem2_145_17, p_wishbone_bd_ram_mem2_145_18,
         p_wishbone_bd_ram_mem2_145_19, p_wishbone_bd_ram_mem2_145_20,
         p_wishbone_bd_ram_mem2_145_21, p_wishbone_bd_ram_mem2_145_22,
         p_wishbone_bd_ram_mem2_145_23, p_wishbone_bd_ram_mem2_146_16,
         p_wishbone_bd_ram_mem2_146_17, p_wishbone_bd_ram_mem2_146_18,
         p_wishbone_bd_ram_mem2_146_19, p_wishbone_bd_ram_mem2_146_20,
         p_wishbone_bd_ram_mem2_146_21, p_wishbone_bd_ram_mem2_146_22,
         p_wishbone_bd_ram_mem2_146_23, p_wishbone_bd_ram_mem2_147_16,
         p_wishbone_bd_ram_mem2_147_17, p_wishbone_bd_ram_mem2_147_18,
         p_wishbone_bd_ram_mem2_147_19, p_wishbone_bd_ram_mem2_147_20,
         p_wishbone_bd_ram_mem2_147_21, p_wishbone_bd_ram_mem2_147_22,
         p_wishbone_bd_ram_mem2_147_23, p_wishbone_bd_ram_mem2_148_16,
         p_wishbone_bd_ram_mem2_148_17, p_wishbone_bd_ram_mem2_148_18,
         p_wishbone_bd_ram_mem2_148_19, p_wishbone_bd_ram_mem2_148_20,
         p_wishbone_bd_ram_mem2_148_21, p_wishbone_bd_ram_mem2_148_22,
         p_wishbone_bd_ram_mem2_148_23, p_wishbone_bd_ram_mem2_149_16,
         p_wishbone_bd_ram_mem2_149_17, p_wishbone_bd_ram_mem2_149_18,
         p_wishbone_bd_ram_mem2_149_19, p_wishbone_bd_ram_mem2_149_20,
         p_wishbone_bd_ram_mem2_149_21, p_wishbone_bd_ram_mem2_149_22,
         p_wishbone_bd_ram_mem2_149_23, p_wishbone_bd_ram_mem2_150_16,
         p_wishbone_bd_ram_mem2_150_17, p_wishbone_bd_ram_mem2_150_18,
         p_wishbone_bd_ram_mem2_150_19, p_wishbone_bd_ram_mem2_150_20,
         p_wishbone_bd_ram_mem2_150_21, p_wishbone_bd_ram_mem2_150_22,
         p_wishbone_bd_ram_mem2_150_23, p_wishbone_bd_ram_mem2_151_16,
         p_wishbone_bd_ram_mem2_151_17, p_wishbone_bd_ram_mem2_151_18,
         p_wishbone_bd_ram_mem2_151_19, p_wishbone_bd_ram_mem2_151_20,
         p_wishbone_bd_ram_mem2_151_21, p_wishbone_bd_ram_mem2_151_22,
         p_wishbone_bd_ram_mem2_151_23, p_wishbone_bd_ram_mem2_152_16,
         p_wishbone_bd_ram_mem2_152_17, p_wishbone_bd_ram_mem2_152_18,
         p_wishbone_bd_ram_mem2_152_19, p_wishbone_bd_ram_mem2_152_20,
         p_wishbone_bd_ram_mem2_152_21, p_wishbone_bd_ram_mem2_152_22,
         p_wishbone_bd_ram_mem2_152_23, p_wishbone_bd_ram_mem2_153_16,
         p_wishbone_bd_ram_mem2_153_17, p_wishbone_bd_ram_mem2_153_18,
         p_wishbone_bd_ram_mem2_153_19, p_wishbone_bd_ram_mem2_153_20,
         p_wishbone_bd_ram_mem2_153_21, p_wishbone_bd_ram_mem2_153_22,
         p_wishbone_bd_ram_mem2_153_23, p_wishbone_bd_ram_mem2_154_16,
         p_wishbone_bd_ram_mem2_154_17, p_wishbone_bd_ram_mem2_154_18,
         p_wishbone_bd_ram_mem2_154_19, p_wishbone_bd_ram_mem2_154_20,
         p_wishbone_bd_ram_mem2_154_21, p_wishbone_bd_ram_mem2_154_22,
         p_wishbone_bd_ram_mem2_154_23, p_wishbone_bd_ram_mem2_155_16,
         p_wishbone_bd_ram_mem2_155_17, p_wishbone_bd_ram_mem2_155_18,
         p_wishbone_bd_ram_mem2_155_19, p_wishbone_bd_ram_mem2_155_20,
         p_wishbone_bd_ram_mem2_155_21, p_wishbone_bd_ram_mem2_155_22,
         p_wishbone_bd_ram_mem2_155_23, p_wishbone_bd_ram_mem2_156_16,
         p_wishbone_bd_ram_mem2_156_17, p_wishbone_bd_ram_mem2_156_18,
         p_wishbone_bd_ram_mem2_156_19, p_wishbone_bd_ram_mem2_156_20,
         p_wishbone_bd_ram_mem2_156_21, p_wishbone_bd_ram_mem2_156_22,
         p_wishbone_bd_ram_mem2_156_23, p_wishbone_bd_ram_mem2_157_16,
         p_wishbone_bd_ram_mem2_157_17, p_wishbone_bd_ram_mem2_157_18,
         p_wishbone_bd_ram_mem2_157_19, p_wishbone_bd_ram_mem2_157_20,
         p_wishbone_bd_ram_mem2_157_21, p_wishbone_bd_ram_mem2_157_22,
         p_wishbone_bd_ram_mem2_157_23, p_wishbone_bd_ram_mem2_158_16,
         p_wishbone_bd_ram_mem2_158_17, p_wishbone_bd_ram_mem2_158_18,
         p_wishbone_bd_ram_mem2_158_19, p_wishbone_bd_ram_mem2_158_20,
         p_wishbone_bd_ram_mem2_158_21, p_wishbone_bd_ram_mem2_158_22,
         p_wishbone_bd_ram_mem2_158_23, p_wishbone_bd_ram_mem2_159_16,
         p_wishbone_bd_ram_mem2_159_17, p_wishbone_bd_ram_mem2_159_18,
         p_wishbone_bd_ram_mem2_159_19, p_wishbone_bd_ram_mem2_159_20,
         p_wishbone_bd_ram_mem2_159_21, p_wishbone_bd_ram_mem2_159_22,
         p_wishbone_bd_ram_mem2_159_23, p_wishbone_bd_ram_mem2_160_16,
         p_wishbone_bd_ram_mem2_160_17, p_wishbone_bd_ram_mem2_160_18,
         p_wishbone_bd_ram_mem2_160_19, p_wishbone_bd_ram_mem2_160_20,
         p_wishbone_bd_ram_mem2_160_21, p_wishbone_bd_ram_mem2_160_22,
         p_wishbone_bd_ram_mem2_160_23, p_wishbone_bd_ram_mem2_161_16,
         p_wishbone_bd_ram_mem2_161_17, p_wishbone_bd_ram_mem2_161_18,
         p_wishbone_bd_ram_mem2_161_19, p_wishbone_bd_ram_mem2_161_20,
         p_wishbone_bd_ram_mem2_161_21, p_wishbone_bd_ram_mem2_161_22,
         p_wishbone_bd_ram_mem2_161_23, p_wishbone_bd_ram_mem2_162_16,
         p_wishbone_bd_ram_mem2_162_17, p_wishbone_bd_ram_mem2_162_18,
         p_wishbone_bd_ram_mem2_162_19, p_wishbone_bd_ram_mem2_162_20,
         p_wishbone_bd_ram_mem2_162_21, p_wishbone_bd_ram_mem2_162_22,
         p_wishbone_bd_ram_mem2_162_23, p_wishbone_bd_ram_mem2_163_16,
         p_wishbone_bd_ram_mem2_163_17, p_wishbone_bd_ram_mem2_163_18,
         p_wishbone_bd_ram_mem2_163_19, p_wishbone_bd_ram_mem2_163_20,
         p_wishbone_bd_ram_mem2_163_21, p_wishbone_bd_ram_mem2_163_22,
         p_wishbone_bd_ram_mem2_163_23, p_wishbone_bd_ram_mem2_164_16,
         p_wishbone_bd_ram_mem2_164_17, p_wishbone_bd_ram_mem2_164_18,
         p_wishbone_bd_ram_mem2_164_19, p_wishbone_bd_ram_mem2_164_20,
         p_wishbone_bd_ram_mem2_164_21, p_wishbone_bd_ram_mem2_164_22,
         p_wishbone_bd_ram_mem2_164_23, p_wishbone_bd_ram_mem2_165_16,
         p_wishbone_bd_ram_mem2_165_17, p_wishbone_bd_ram_mem2_165_18,
         p_wishbone_bd_ram_mem2_165_19, p_wishbone_bd_ram_mem2_165_20,
         p_wishbone_bd_ram_mem2_165_21, p_wishbone_bd_ram_mem2_165_22,
         p_wishbone_bd_ram_mem2_165_23, p_wishbone_bd_ram_mem2_166_16,
         p_wishbone_bd_ram_mem2_166_17, p_wishbone_bd_ram_mem2_166_18,
         p_wishbone_bd_ram_mem2_166_19, p_wishbone_bd_ram_mem2_166_20,
         p_wishbone_bd_ram_mem2_166_21, p_wishbone_bd_ram_mem2_166_22,
         p_wishbone_bd_ram_mem2_166_23, p_wishbone_bd_ram_mem2_167_16,
         p_wishbone_bd_ram_mem2_167_17, p_wishbone_bd_ram_mem2_167_18,
         p_wishbone_bd_ram_mem2_167_19, p_wishbone_bd_ram_mem2_167_20,
         p_wishbone_bd_ram_mem2_167_21, p_wishbone_bd_ram_mem2_167_22,
         p_wishbone_bd_ram_mem2_167_23, p_wishbone_bd_ram_mem2_168_16,
         p_wishbone_bd_ram_mem2_168_17, p_wishbone_bd_ram_mem2_168_18,
         p_wishbone_bd_ram_mem2_168_19, p_wishbone_bd_ram_mem2_168_20,
         p_wishbone_bd_ram_mem2_168_21, p_wishbone_bd_ram_mem2_168_22,
         p_wishbone_bd_ram_mem2_168_23, p_wishbone_bd_ram_mem2_169_16,
         p_wishbone_bd_ram_mem2_169_17, p_wishbone_bd_ram_mem2_169_18,
         p_wishbone_bd_ram_mem2_169_19, p_wishbone_bd_ram_mem2_169_20,
         p_wishbone_bd_ram_mem2_169_21, p_wishbone_bd_ram_mem2_169_22,
         p_wishbone_bd_ram_mem2_169_23, p_wishbone_bd_ram_mem2_170_16,
         p_wishbone_bd_ram_mem2_170_17, p_wishbone_bd_ram_mem2_170_18,
         p_wishbone_bd_ram_mem2_170_19, p_wishbone_bd_ram_mem2_170_20,
         p_wishbone_bd_ram_mem2_170_21, p_wishbone_bd_ram_mem2_170_22,
         p_wishbone_bd_ram_mem2_170_23, p_wishbone_bd_ram_mem2_171_16,
         p_wishbone_bd_ram_mem2_171_17, p_wishbone_bd_ram_mem2_171_18,
         p_wishbone_bd_ram_mem2_171_19, p_wishbone_bd_ram_mem2_171_20,
         p_wishbone_bd_ram_mem2_171_21, p_wishbone_bd_ram_mem2_171_22,
         p_wishbone_bd_ram_mem2_171_23, p_wishbone_bd_ram_mem2_172_16,
         p_wishbone_bd_ram_mem2_172_17, p_wishbone_bd_ram_mem2_172_18,
         p_wishbone_bd_ram_mem2_172_19, p_wishbone_bd_ram_mem2_172_20,
         p_wishbone_bd_ram_mem2_172_21, p_wishbone_bd_ram_mem2_172_22,
         p_wishbone_bd_ram_mem2_172_23, p_wishbone_bd_ram_mem2_173_16,
         p_wishbone_bd_ram_mem2_173_17, p_wishbone_bd_ram_mem2_173_18,
         p_wishbone_bd_ram_mem2_173_19, p_wishbone_bd_ram_mem2_173_20,
         p_wishbone_bd_ram_mem2_173_21, p_wishbone_bd_ram_mem2_173_22,
         p_wishbone_bd_ram_mem2_173_23, p_wishbone_bd_ram_mem2_174_16,
         p_wishbone_bd_ram_mem2_174_17, p_wishbone_bd_ram_mem2_174_18,
         p_wishbone_bd_ram_mem2_174_19, p_wishbone_bd_ram_mem2_174_20,
         p_wishbone_bd_ram_mem2_174_21, p_wishbone_bd_ram_mem2_174_22,
         p_wishbone_bd_ram_mem2_174_23, p_wishbone_bd_ram_mem2_175_16,
         p_wishbone_bd_ram_mem2_175_17, p_wishbone_bd_ram_mem2_175_18,
         p_wishbone_bd_ram_mem2_175_19, p_wishbone_bd_ram_mem2_175_20,
         p_wishbone_bd_ram_mem2_175_21, p_wishbone_bd_ram_mem2_175_22,
         p_wishbone_bd_ram_mem2_175_23, p_wishbone_bd_ram_mem2_176_16,
         p_wishbone_bd_ram_mem2_176_17, p_wishbone_bd_ram_mem2_176_18,
         p_wishbone_bd_ram_mem2_176_19, p_wishbone_bd_ram_mem2_176_20,
         p_wishbone_bd_ram_mem2_176_21, p_wishbone_bd_ram_mem2_176_22,
         p_wishbone_bd_ram_mem2_176_23, p_wishbone_bd_ram_mem2_177_16,
         p_wishbone_bd_ram_mem2_177_17, p_wishbone_bd_ram_mem2_177_18,
         p_wishbone_bd_ram_mem2_177_19, p_wishbone_bd_ram_mem2_177_20,
         p_wishbone_bd_ram_mem2_177_21, p_wishbone_bd_ram_mem2_177_22,
         p_wishbone_bd_ram_mem2_177_23, p_wishbone_bd_ram_mem2_178_16,
         p_wishbone_bd_ram_mem2_178_17, p_wishbone_bd_ram_mem2_178_18,
         p_wishbone_bd_ram_mem2_178_19, p_wishbone_bd_ram_mem2_178_20,
         p_wishbone_bd_ram_mem2_178_21, p_wishbone_bd_ram_mem2_178_22,
         p_wishbone_bd_ram_mem2_178_23, p_wishbone_bd_ram_mem2_179_16,
         p_wishbone_bd_ram_mem2_179_17, p_wishbone_bd_ram_mem2_179_18,
         p_wishbone_bd_ram_mem2_179_19, p_wishbone_bd_ram_mem2_179_20,
         p_wishbone_bd_ram_mem2_179_21, p_wishbone_bd_ram_mem2_179_22,
         p_wishbone_bd_ram_mem2_179_23, p_wishbone_bd_ram_mem2_180_16,
         p_wishbone_bd_ram_mem2_180_17, p_wishbone_bd_ram_mem2_180_18,
         p_wishbone_bd_ram_mem2_180_19, p_wishbone_bd_ram_mem2_180_20,
         p_wishbone_bd_ram_mem2_180_21, p_wishbone_bd_ram_mem2_180_22,
         p_wishbone_bd_ram_mem2_180_23, p_wishbone_bd_ram_mem2_181_16,
         p_wishbone_bd_ram_mem2_181_17, p_wishbone_bd_ram_mem2_181_18,
         p_wishbone_bd_ram_mem2_181_19, p_wishbone_bd_ram_mem2_181_20,
         p_wishbone_bd_ram_mem2_181_21, p_wishbone_bd_ram_mem2_181_22,
         p_wishbone_bd_ram_mem2_181_23, p_wishbone_bd_ram_mem2_182_16,
         p_wishbone_bd_ram_mem2_182_17, p_wishbone_bd_ram_mem2_182_18,
         p_wishbone_bd_ram_mem2_182_19, p_wishbone_bd_ram_mem2_182_20,
         p_wishbone_bd_ram_mem2_182_21, p_wishbone_bd_ram_mem2_182_22,
         p_wishbone_bd_ram_mem2_182_23, p_wishbone_bd_ram_mem2_183_16,
         p_wishbone_bd_ram_mem2_183_17, p_wishbone_bd_ram_mem2_183_18,
         p_wishbone_bd_ram_mem2_183_19, p_wishbone_bd_ram_mem2_183_20,
         p_wishbone_bd_ram_mem2_183_21, p_wishbone_bd_ram_mem2_183_22,
         p_wishbone_bd_ram_mem2_183_23, p_wishbone_bd_ram_mem2_184_16,
         p_wishbone_bd_ram_mem2_184_17, p_wishbone_bd_ram_mem2_184_18,
         p_wishbone_bd_ram_mem2_184_19, p_wishbone_bd_ram_mem2_184_20,
         p_wishbone_bd_ram_mem2_184_21, p_wishbone_bd_ram_mem2_184_22,
         p_wishbone_bd_ram_mem2_184_23, p_wishbone_bd_ram_mem2_185_16,
         p_wishbone_bd_ram_mem2_185_17, p_wishbone_bd_ram_mem2_185_18,
         p_wishbone_bd_ram_mem2_185_19, p_wishbone_bd_ram_mem2_185_20,
         p_wishbone_bd_ram_mem2_185_21, p_wishbone_bd_ram_mem2_185_22,
         p_wishbone_bd_ram_mem2_185_23, p_wishbone_bd_ram_mem2_186_16,
         p_wishbone_bd_ram_mem2_186_17, p_wishbone_bd_ram_mem2_186_18,
         p_wishbone_bd_ram_mem2_186_19, p_wishbone_bd_ram_mem2_186_20,
         p_wishbone_bd_ram_mem2_186_21, p_wishbone_bd_ram_mem2_186_22,
         p_wishbone_bd_ram_mem2_186_23, p_wishbone_bd_ram_mem2_187_16,
         p_wishbone_bd_ram_mem2_187_17, p_wishbone_bd_ram_mem2_187_18,
         p_wishbone_bd_ram_mem2_187_19, p_wishbone_bd_ram_mem2_187_20,
         p_wishbone_bd_ram_mem2_187_21, p_wishbone_bd_ram_mem2_187_22,
         p_wishbone_bd_ram_mem2_187_23, p_wishbone_bd_ram_mem2_188_16,
         p_wishbone_bd_ram_mem2_188_17, p_wishbone_bd_ram_mem2_188_18,
         p_wishbone_bd_ram_mem2_188_19, p_wishbone_bd_ram_mem2_188_20,
         p_wishbone_bd_ram_mem2_188_21, p_wishbone_bd_ram_mem2_188_22,
         p_wishbone_bd_ram_mem2_188_23, p_wishbone_bd_ram_mem2_189_16,
         p_wishbone_bd_ram_mem2_189_17, p_wishbone_bd_ram_mem2_189_18,
         p_wishbone_bd_ram_mem2_189_19, p_wishbone_bd_ram_mem2_189_20,
         p_wishbone_bd_ram_mem2_189_21, p_wishbone_bd_ram_mem2_189_22,
         p_wishbone_bd_ram_mem2_189_23, p_wishbone_bd_ram_mem2_190_16,
         p_wishbone_bd_ram_mem2_190_17, p_wishbone_bd_ram_mem2_190_18,
         p_wishbone_bd_ram_mem2_190_19, p_wishbone_bd_ram_mem2_190_20,
         p_wishbone_bd_ram_mem2_190_21, p_wishbone_bd_ram_mem2_190_22,
         p_wishbone_bd_ram_mem2_190_23, p_wishbone_bd_ram_mem2_191_16,
         p_wishbone_bd_ram_mem2_191_17, p_wishbone_bd_ram_mem2_191_18,
         p_wishbone_bd_ram_mem2_191_19, p_wishbone_bd_ram_mem2_191_20,
         p_wishbone_bd_ram_mem2_191_21, p_wishbone_bd_ram_mem2_191_22,
         p_wishbone_bd_ram_mem2_191_23, p_wishbone_bd_ram_mem2_192_16,
         p_wishbone_bd_ram_mem2_192_17, p_wishbone_bd_ram_mem2_192_18,
         p_wishbone_bd_ram_mem2_192_19, p_wishbone_bd_ram_mem2_192_20,
         p_wishbone_bd_ram_mem2_192_21, p_wishbone_bd_ram_mem2_192_22,
         p_wishbone_bd_ram_mem2_192_23, p_wishbone_bd_ram_mem2_193_16,
         p_wishbone_bd_ram_mem2_193_17, p_wishbone_bd_ram_mem2_193_18,
         p_wishbone_bd_ram_mem2_193_19, p_wishbone_bd_ram_mem2_193_20,
         p_wishbone_bd_ram_mem2_193_21, p_wishbone_bd_ram_mem2_193_22,
         p_wishbone_bd_ram_mem2_193_23, p_wishbone_bd_ram_mem2_194_16,
         p_wishbone_bd_ram_mem2_194_17, p_wishbone_bd_ram_mem2_194_18,
         p_wishbone_bd_ram_mem2_194_19, p_wishbone_bd_ram_mem2_194_20,
         p_wishbone_bd_ram_mem2_194_21, p_wishbone_bd_ram_mem2_194_22,
         p_wishbone_bd_ram_mem2_194_23, p_wishbone_bd_ram_mem2_195_16,
         p_wishbone_bd_ram_mem2_195_17, p_wishbone_bd_ram_mem2_195_18,
         p_wishbone_bd_ram_mem2_195_19, p_wishbone_bd_ram_mem2_195_20,
         p_wishbone_bd_ram_mem2_195_21, p_wishbone_bd_ram_mem2_195_22,
         p_wishbone_bd_ram_mem2_195_23, p_wishbone_bd_ram_mem2_196_16,
         p_wishbone_bd_ram_mem2_196_17, p_wishbone_bd_ram_mem2_196_18,
         p_wishbone_bd_ram_mem2_196_19, p_wishbone_bd_ram_mem2_196_20,
         p_wishbone_bd_ram_mem2_196_21, p_wishbone_bd_ram_mem2_196_22,
         p_wishbone_bd_ram_mem2_196_23, p_wishbone_bd_ram_mem2_197_16,
         p_wishbone_bd_ram_mem2_197_17, p_wishbone_bd_ram_mem2_197_18,
         p_wishbone_bd_ram_mem2_197_19, p_wishbone_bd_ram_mem2_197_20,
         p_wishbone_bd_ram_mem2_197_21, p_wishbone_bd_ram_mem2_197_22,
         p_wishbone_bd_ram_mem2_197_23, p_wishbone_bd_ram_mem2_198_16,
         p_wishbone_bd_ram_mem2_198_17, p_wishbone_bd_ram_mem2_198_18,
         p_wishbone_bd_ram_mem2_198_19, p_wishbone_bd_ram_mem2_198_20,
         p_wishbone_bd_ram_mem2_198_21, p_wishbone_bd_ram_mem2_198_22,
         p_wishbone_bd_ram_mem2_198_23, p_wishbone_bd_ram_mem2_199_16,
         p_wishbone_bd_ram_mem2_199_17, p_wishbone_bd_ram_mem2_199_18,
         p_wishbone_bd_ram_mem2_199_19, p_wishbone_bd_ram_mem2_199_20,
         p_wishbone_bd_ram_mem2_199_21, p_wishbone_bd_ram_mem2_199_22,
         p_wishbone_bd_ram_mem2_199_23, p_wishbone_bd_ram_mem2_200_16,
         p_wishbone_bd_ram_mem2_200_17, p_wishbone_bd_ram_mem2_200_18,
         p_wishbone_bd_ram_mem2_200_19, p_wishbone_bd_ram_mem2_200_20,
         p_wishbone_bd_ram_mem2_200_21, p_wishbone_bd_ram_mem2_200_22,
         p_wishbone_bd_ram_mem2_200_23, p_wishbone_bd_ram_mem2_201_16,
         p_wishbone_bd_ram_mem2_201_17, p_wishbone_bd_ram_mem2_201_18,
         p_wishbone_bd_ram_mem2_201_19, p_wishbone_bd_ram_mem2_201_20,
         p_wishbone_bd_ram_mem2_201_21, p_wishbone_bd_ram_mem2_201_22,
         p_wishbone_bd_ram_mem2_201_23, p_wishbone_bd_ram_mem2_202_16,
         p_wishbone_bd_ram_mem2_202_17, p_wishbone_bd_ram_mem2_202_18,
         p_wishbone_bd_ram_mem2_202_19, p_wishbone_bd_ram_mem2_202_20,
         p_wishbone_bd_ram_mem2_202_21, p_wishbone_bd_ram_mem2_202_22,
         p_wishbone_bd_ram_mem2_202_23, p_wishbone_bd_ram_mem2_203_16,
         p_wishbone_bd_ram_mem2_203_17, p_wishbone_bd_ram_mem2_203_18,
         p_wishbone_bd_ram_mem2_203_19, p_wishbone_bd_ram_mem2_203_20,
         p_wishbone_bd_ram_mem2_203_21, p_wishbone_bd_ram_mem2_203_22,
         p_wishbone_bd_ram_mem2_203_23, p_wishbone_bd_ram_mem2_204_16,
         p_wishbone_bd_ram_mem2_204_17, p_wishbone_bd_ram_mem2_204_18,
         p_wishbone_bd_ram_mem2_204_19, p_wishbone_bd_ram_mem2_204_20,
         p_wishbone_bd_ram_mem2_204_21, p_wishbone_bd_ram_mem2_204_22,
         p_wishbone_bd_ram_mem2_204_23, p_wishbone_bd_ram_mem2_205_16,
         p_wishbone_bd_ram_mem2_205_17, p_wishbone_bd_ram_mem2_205_18,
         p_wishbone_bd_ram_mem2_205_19, p_wishbone_bd_ram_mem2_205_20,
         p_wishbone_bd_ram_mem2_205_21, p_wishbone_bd_ram_mem2_205_22,
         p_wishbone_bd_ram_mem2_205_23, p_wishbone_bd_ram_mem2_206_16,
         p_wishbone_bd_ram_mem2_206_17, p_wishbone_bd_ram_mem2_206_18,
         p_wishbone_bd_ram_mem2_206_19, p_wishbone_bd_ram_mem2_206_20,
         p_wishbone_bd_ram_mem2_206_21, p_wishbone_bd_ram_mem2_206_22,
         p_wishbone_bd_ram_mem2_206_23, p_wishbone_bd_ram_mem2_207_16,
         p_wishbone_bd_ram_mem2_207_17, p_wishbone_bd_ram_mem2_207_18,
         p_wishbone_bd_ram_mem2_207_19, p_wishbone_bd_ram_mem2_207_20,
         p_wishbone_bd_ram_mem2_207_21, p_wishbone_bd_ram_mem2_207_22,
         p_wishbone_bd_ram_mem2_207_23, p_wishbone_bd_ram_mem2_208_16,
         p_wishbone_bd_ram_mem2_208_17, p_wishbone_bd_ram_mem2_208_18,
         p_wishbone_bd_ram_mem2_208_19, p_wishbone_bd_ram_mem2_208_20,
         p_wishbone_bd_ram_mem2_208_21, p_wishbone_bd_ram_mem2_208_22,
         p_wishbone_bd_ram_mem2_208_23, p_wishbone_bd_ram_mem2_209_16,
         p_wishbone_bd_ram_mem2_209_17, p_wishbone_bd_ram_mem2_209_18,
         p_wishbone_bd_ram_mem2_209_19, p_wishbone_bd_ram_mem2_209_20,
         p_wishbone_bd_ram_mem2_209_21, p_wishbone_bd_ram_mem2_209_22,
         p_wishbone_bd_ram_mem2_209_23, p_wishbone_bd_ram_mem2_210_16,
         p_wishbone_bd_ram_mem2_210_17, p_wishbone_bd_ram_mem2_210_18,
         p_wishbone_bd_ram_mem2_210_19, p_wishbone_bd_ram_mem2_210_20,
         p_wishbone_bd_ram_mem2_210_21, p_wishbone_bd_ram_mem2_210_22,
         p_wishbone_bd_ram_mem2_210_23, p_wishbone_bd_ram_mem2_211_16,
         p_wishbone_bd_ram_mem2_211_17, p_wishbone_bd_ram_mem2_211_18,
         p_wishbone_bd_ram_mem2_211_19, p_wishbone_bd_ram_mem2_211_20,
         p_wishbone_bd_ram_mem2_211_21, p_wishbone_bd_ram_mem2_211_22,
         p_wishbone_bd_ram_mem2_211_23, p_wishbone_bd_ram_mem2_212_16,
         p_wishbone_bd_ram_mem2_212_17, p_wishbone_bd_ram_mem2_212_18,
         p_wishbone_bd_ram_mem2_212_19, p_wishbone_bd_ram_mem2_212_20,
         p_wishbone_bd_ram_mem2_212_21, p_wishbone_bd_ram_mem2_212_22,
         p_wishbone_bd_ram_mem2_212_23, p_wishbone_bd_ram_mem2_213_16,
         p_wishbone_bd_ram_mem2_213_17, p_wishbone_bd_ram_mem2_213_18,
         p_wishbone_bd_ram_mem2_213_19, p_wishbone_bd_ram_mem2_213_20,
         p_wishbone_bd_ram_mem2_213_21, p_wishbone_bd_ram_mem2_213_22,
         p_wishbone_bd_ram_mem2_213_23, p_wishbone_bd_ram_mem2_214_16,
         p_wishbone_bd_ram_mem2_214_17, p_wishbone_bd_ram_mem2_214_18,
         p_wishbone_bd_ram_mem2_214_19, p_wishbone_bd_ram_mem2_214_20,
         p_wishbone_bd_ram_mem2_214_21, p_wishbone_bd_ram_mem2_214_22,
         p_wishbone_bd_ram_mem2_214_23, p_wishbone_bd_ram_mem2_215_16,
         p_wishbone_bd_ram_mem2_215_17, p_wishbone_bd_ram_mem2_215_18,
         p_wishbone_bd_ram_mem2_215_19, p_wishbone_bd_ram_mem2_215_20,
         p_wishbone_bd_ram_mem2_215_21, p_wishbone_bd_ram_mem2_215_22,
         p_wishbone_bd_ram_mem2_215_23, p_wishbone_bd_ram_mem2_216_16,
         p_wishbone_bd_ram_mem2_216_17, p_wishbone_bd_ram_mem2_216_18,
         p_wishbone_bd_ram_mem2_216_19, p_wishbone_bd_ram_mem2_216_20,
         p_wishbone_bd_ram_mem2_216_21, p_wishbone_bd_ram_mem2_216_22,
         p_wishbone_bd_ram_mem2_216_23, p_wishbone_bd_ram_mem2_217_16,
         p_wishbone_bd_ram_mem2_217_17, p_wishbone_bd_ram_mem2_217_18,
         p_wishbone_bd_ram_mem2_217_19, p_wishbone_bd_ram_mem2_217_20,
         p_wishbone_bd_ram_mem2_217_21, p_wishbone_bd_ram_mem2_217_22,
         p_wishbone_bd_ram_mem2_217_23, p_wishbone_bd_ram_mem2_218_16,
         p_wishbone_bd_ram_mem2_218_17, p_wishbone_bd_ram_mem2_218_18,
         p_wishbone_bd_ram_mem2_218_19, p_wishbone_bd_ram_mem2_218_20,
         p_wishbone_bd_ram_mem2_218_21, p_wishbone_bd_ram_mem2_218_22,
         p_wishbone_bd_ram_mem2_218_23, p_wishbone_bd_ram_mem2_219_16,
         p_wishbone_bd_ram_mem2_219_17, p_wishbone_bd_ram_mem2_219_18,
         p_wishbone_bd_ram_mem2_219_19, p_wishbone_bd_ram_mem2_219_20,
         p_wishbone_bd_ram_mem2_219_21, p_wishbone_bd_ram_mem2_219_22,
         p_wishbone_bd_ram_mem2_219_23, p_wishbone_bd_ram_mem2_220_16,
         p_wishbone_bd_ram_mem2_220_17, p_wishbone_bd_ram_mem2_220_18,
         p_wishbone_bd_ram_mem2_220_19, p_wishbone_bd_ram_mem2_220_20,
         p_wishbone_bd_ram_mem2_220_21, p_wishbone_bd_ram_mem2_220_22,
         p_wishbone_bd_ram_mem2_220_23, p_wishbone_bd_ram_mem2_221_16,
         p_wishbone_bd_ram_mem2_221_17, p_wishbone_bd_ram_mem2_221_18,
         p_wishbone_bd_ram_mem2_221_19, p_wishbone_bd_ram_mem2_221_20,
         p_wishbone_bd_ram_mem2_221_21, p_wishbone_bd_ram_mem2_221_22,
         p_wishbone_bd_ram_mem2_221_23, p_wishbone_bd_ram_mem2_222_16,
         p_wishbone_bd_ram_mem2_222_17, p_wishbone_bd_ram_mem2_222_18,
         p_wishbone_bd_ram_mem2_222_19, p_wishbone_bd_ram_mem2_222_20,
         p_wishbone_bd_ram_mem2_222_21, p_wishbone_bd_ram_mem2_222_22,
         p_wishbone_bd_ram_mem2_222_23, p_wishbone_bd_ram_mem2_223_16,
         p_wishbone_bd_ram_mem2_223_17, p_wishbone_bd_ram_mem2_223_18,
         p_wishbone_bd_ram_mem2_223_19, p_wishbone_bd_ram_mem2_223_20,
         p_wishbone_bd_ram_mem2_223_21, p_wishbone_bd_ram_mem2_223_22,
         p_wishbone_bd_ram_mem2_223_23, p_wishbone_bd_ram_mem2_224_16,
         p_wishbone_bd_ram_mem2_224_17, p_wishbone_bd_ram_mem2_224_18,
         p_wishbone_bd_ram_mem2_224_19, p_wishbone_bd_ram_mem2_224_20,
         p_wishbone_bd_ram_mem2_224_21, p_wishbone_bd_ram_mem2_224_22,
         p_wishbone_bd_ram_mem2_224_23, p_wishbone_bd_ram_mem2_225_16,
         p_wishbone_bd_ram_mem2_225_17, p_wishbone_bd_ram_mem2_225_18,
         p_wishbone_bd_ram_mem2_225_19, p_wishbone_bd_ram_mem2_225_20,
         p_wishbone_bd_ram_mem2_225_21, p_wishbone_bd_ram_mem2_225_22,
         p_wishbone_bd_ram_mem2_225_23, p_wishbone_bd_ram_mem2_226_16,
         p_wishbone_bd_ram_mem2_226_17, p_wishbone_bd_ram_mem2_226_18,
         p_wishbone_bd_ram_mem2_226_19, p_wishbone_bd_ram_mem2_226_20,
         p_wishbone_bd_ram_mem2_226_21, p_wishbone_bd_ram_mem2_226_22,
         p_wishbone_bd_ram_mem2_226_23, p_wishbone_bd_ram_mem2_227_16,
         p_wishbone_bd_ram_mem2_227_17, p_wishbone_bd_ram_mem2_227_18,
         p_wishbone_bd_ram_mem2_227_19, p_wishbone_bd_ram_mem2_227_20,
         p_wishbone_bd_ram_mem2_227_21, p_wishbone_bd_ram_mem2_227_22,
         p_wishbone_bd_ram_mem2_227_23, p_wishbone_bd_ram_mem2_228_16,
         p_wishbone_bd_ram_mem2_228_17, p_wishbone_bd_ram_mem2_228_18,
         p_wishbone_bd_ram_mem2_228_19, p_wishbone_bd_ram_mem2_228_20,
         p_wishbone_bd_ram_mem2_228_21, p_wishbone_bd_ram_mem2_228_22,
         p_wishbone_bd_ram_mem2_228_23, p_wishbone_bd_ram_mem2_229_16,
         p_wishbone_bd_ram_mem2_229_17, p_wishbone_bd_ram_mem2_229_18,
         p_wishbone_bd_ram_mem2_229_19, p_wishbone_bd_ram_mem2_229_20,
         p_wishbone_bd_ram_mem2_229_21, p_wishbone_bd_ram_mem2_229_22,
         p_wishbone_bd_ram_mem2_229_23, p_wishbone_bd_ram_mem2_230_16,
         p_wishbone_bd_ram_mem2_230_17, p_wishbone_bd_ram_mem2_230_18,
         p_wishbone_bd_ram_mem2_230_19, p_wishbone_bd_ram_mem2_230_20,
         p_wishbone_bd_ram_mem2_230_21, p_wishbone_bd_ram_mem2_230_22,
         p_wishbone_bd_ram_mem2_230_23, p_wishbone_bd_ram_mem2_231_16,
         p_wishbone_bd_ram_mem2_231_17, p_wishbone_bd_ram_mem2_231_18,
         p_wishbone_bd_ram_mem2_231_19, p_wishbone_bd_ram_mem2_231_20,
         p_wishbone_bd_ram_mem2_231_21, p_wishbone_bd_ram_mem2_231_22,
         p_wishbone_bd_ram_mem2_231_23, p_wishbone_bd_ram_mem2_232_16,
         p_wishbone_bd_ram_mem2_232_17, p_wishbone_bd_ram_mem2_232_18,
         p_wishbone_bd_ram_mem2_232_19, p_wishbone_bd_ram_mem2_232_20,
         p_wishbone_bd_ram_mem2_232_21, p_wishbone_bd_ram_mem2_232_22,
         p_wishbone_bd_ram_mem2_232_23, p_wishbone_bd_ram_mem2_233_16,
         p_wishbone_bd_ram_mem2_233_17, p_wishbone_bd_ram_mem2_233_18,
         p_wishbone_bd_ram_mem2_233_19, p_wishbone_bd_ram_mem2_233_20,
         p_wishbone_bd_ram_mem2_233_21, p_wishbone_bd_ram_mem2_233_22,
         p_wishbone_bd_ram_mem2_233_23, p_wishbone_bd_ram_mem2_234_16,
         p_wishbone_bd_ram_mem2_234_17, p_wishbone_bd_ram_mem2_234_18,
         p_wishbone_bd_ram_mem2_234_19, p_wishbone_bd_ram_mem2_234_20,
         p_wishbone_bd_ram_mem2_234_21, p_wishbone_bd_ram_mem2_234_22,
         p_wishbone_bd_ram_mem2_234_23, p_wishbone_bd_ram_mem2_235_16,
         p_wishbone_bd_ram_mem2_235_17, p_wishbone_bd_ram_mem2_235_18,
         p_wishbone_bd_ram_mem2_235_19, p_wishbone_bd_ram_mem2_235_20,
         p_wishbone_bd_ram_mem2_235_21, p_wishbone_bd_ram_mem2_235_22,
         p_wishbone_bd_ram_mem2_235_23, p_wishbone_bd_ram_mem2_236_16,
         p_wishbone_bd_ram_mem2_236_17, p_wishbone_bd_ram_mem2_236_18,
         p_wishbone_bd_ram_mem2_236_19, p_wishbone_bd_ram_mem2_236_20,
         p_wishbone_bd_ram_mem2_236_21, p_wishbone_bd_ram_mem2_236_22,
         p_wishbone_bd_ram_mem2_236_23, p_wishbone_bd_ram_mem2_237_16,
         p_wishbone_bd_ram_mem2_237_17, p_wishbone_bd_ram_mem2_237_18,
         p_wishbone_bd_ram_mem2_237_19, p_wishbone_bd_ram_mem2_237_20,
         p_wishbone_bd_ram_mem2_237_21, p_wishbone_bd_ram_mem2_237_22,
         p_wishbone_bd_ram_mem2_237_23, p_wishbone_bd_ram_mem2_238_16,
         p_wishbone_bd_ram_mem2_238_17, p_wishbone_bd_ram_mem2_238_18,
         p_wishbone_bd_ram_mem2_238_19, p_wishbone_bd_ram_mem2_238_20,
         p_wishbone_bd_ram_mem2_238_21, p_wishbone_bd_ram_mem2_238_22,
         p_wishbone_bd_ram_mem2_238_23, p_wishbone_bd_ram_mem2_239_16,
         p_wishbone_bd_ram_mem2_239_17, p_wishbone_bd_ram_mem2_239_18,
         p_wishbone_bd_ram_mem2_239_19, p_wishbone_bd_ram_mem2_239_20,
         p_wishbone_bd_ram_mem2_239_21, p_wishbone_bd_ram_mem2_239_22,
         p_wishbone_bd_ram_mem2_239_23, p_wishbone_bd_ram_mem2_240_16,
         p_wishbone_bd_ram_mem2_240_17, p_wishbone_bd_ram_mem2_240_18,
         p_wishbone_bd_ram_mem2_240_19, p_wishbone_bd_ram_mem2_240_20,
         p_wishbone_bd_ram_mem2_240_21, p_wishbone_bd_ram_mem2_240_22,
         p_wishbone_bd_ram_mem2_240_23, p_wishbone_bd_ram_mem2_241_16,
         p_wishbone_bd_ram_mem2_241_17, p_wishbone_bd_ram_mem2_241_18,
         p_wishbone_bd_ram_mem2_241_19, p_wishbone_bd_ram_mem2_241_20,
         p_wishbone_bd_ram_mem2_241_21, p_wishbone_bd_ram_mem2_241_22,
         p_wishbone_bd_ram_mem2_241_23, p_wishbone_bd_ram_mem2_242_16,
         p_wishbone_bd_ram_mem2_242_17, p_wishbone_bd_ram_mem2_242_18,
         p_wishbone_bd_ram_mem2_242_19, p_wishbone_bd_ram_mem2_242_20,
         p_wishbone_bd_ram_mem2_242_21, p_wishbone_bd_ram_mem2_242_22,
         p_wishbone_bd_ram_mem2_242_23, p_wishbone_bd_ram_mem2_243_16,
         p_wishbone_bd_ram_mem2_243_17, p_wishbone_bd_ram_mem2_243_18,
         p_wishbone_bd_ram_mem2_243_19, p_wishbone_bd_ram_mem2_243_20,
         p_wishbone_bd_ram_mem2_243_21, p_wishbone_bd_ram_mem2_243_22,
         p_wishbone_bd_ram_mem2_243_23, p_wishbone_bd_ram_mem2_244_16,
         p_wishbone_bd_ram_mem2_244_17, p_wishbone_bd_ram_mem2_244_18,
         p_wishbone_bd_ram_mem2_244_19, p_wishbone_bd_ram_mem2_244_20,
         p_wishbone_bd_ram_mem2_244_21, p_wishbone_bd_ram_mem2_244_22,
         p_wishbone_bd_ram_mem2_244_23, p_wishbone_bd_ram_mem2_245_16,
         p_wishbone_bd_ram_mem2_245_17, p_wishbone_bd_ram_mem2_245_18,
         p_wishbone_bd_ram_mem2_245_19, p_wishbone_bd_ram_mem2_245_20,
         p_wishbone_bd_ram_mem2_245_21, p_wishbone_bd_ram_mem2_245_22,
         p_wishbone_bd_ram_mem2_245_23, p_wishbone_bd_ram_mem2_246_16,
         p_wishbone_bd_ram_mem2_246_17, p_wishbone_bd_ram_mem2_246_18,
         p_wishbone_bd_ram_mem2_246_19, p_wishbone_bd_ram_mem2_246_20,
         p_wishbone_bd_ram_mem2_246_21, p_wishbone_bd_ram_mem2_246_22,
         p_wishbone_bd_ram_mem2_246_23, p_wishbone_bd_ram_mem2_247_16,
         p_wishbone_bd_ram_mem2_247_17, p_wishbone_bd_ram_mem2_247_18,
         p_wishbone_bd_ram_mem2_247_19, p_wishbone_bd_ram_mem2_247_20,
         p_wishbone_bd_ram_mem2_247_21, p_wishbone_bd_ram_mem2_247_22,
         p_wishbone_bd_ram_mem2_247_23, p_wishbone_bd_ram_mem2_248_16,
         p_wishbone_bd_ram_mem2_248_17, p_wishbone_bd_ram_mem2_248_18,
         p_wishbone_bd_ram_mem2_248_19, p_wishbone_bd_ram_mem2_248_20,
         p_wishbone_bd_ram_mem2_248_21, p_wishbone_bd_ram_mem2_248_22,
         p_wishbone_bd_ram_mem2_248_23, p_wishbone_bd_ram_mem2_249_16,
         p_wishbone_bd_ram_mem2_249_17, p_wishbone_bd_ram_mem2_249_18,
         p_wishbone_bd_ram_mem2_249_19, p_wishbone_bd_ram_mem2_249_20,
         p_wishbone_bd_ram_mem2_249_21, p_wishbone_bd_ram_mem2_249_22,
         p_wishbone_bd_ram_mem2_249_23, p_wishbone_bd_ram_mem2_250_16,
         p_wishbone_bd_ram_mem2_250_17, p_wishbone_bd_ram_mem2_250_18,
         p_wishbone_bd_ram_mem2_250_19, p_wishbone_bd_ram_mem2_250_20,
         p_wishbone_bd_ram_mem2_250_21, p_wishbone_bd_ram_mem2_250_22,
         p_wishbone_bd_ram_mem2_250_23, p_wishbone_bd_ram_mem2_251_16,
         p_wishbone_bd_ram_mem2_251_17, p_wishbone_bd_ram_mem2_251_18,
         p_wishbone_bd_ram_mem2_251_19, p_wishbone_bd_ram_mem2_251_20,
         p_wishbone_bd_ram_mem2_251_21, p_wishbone_bd_ram_mem2_251_22,
         p_wishbone_bd_ram_mem2_251_23, p_wishbone_bd_ram_mem2_252_16,
         p_wishbone_bd_ram_mem2_252_17, p_wishbone_bd_ram_mem2_252_18,
         p_wishbone_bd_ram_mem2_252_19, p_wishbone_bd_ram_mem2_252_20,
         p_wishbone_bd_ram_mem2_252_21, p_wishbone_bd_ram_mem2_252_22,
         p_wishbone_bd_ram_mem2_252_23, p_wishbone_bd_ram_mem2_253_16,
         p_wishbone_bd_ram_mem2_253_17, p_wishbone_bd_ram_mem2_253_18,
         p_wishbone_bd_ram_mem2_253_19, p_wishbone_bd_ram_mem2_253_20,
         p_wishbone_bd_ram_mem2_253_21, p_wishbone_bd_ram_mem2_253_22,
         p_wishbone_bd_ram_mem2_253_23, p_wishbone_bd_ram_mem2_254_16,
         p_wishbone_bd_ram_mem2_254_17, p_wishbone_bd_ram_mem2_254_18,
         p_wishbone_bd_ram_mem2_254_19, p_wishbone_bd_ram_mem2_254_20,
         p_wishbone_bd_ram_mem2_254_21, p_wishbone_bd_ram_mem2_254_22,
         p_wishbone_bd_ram_mem2_254_23, p_wishbone_bd_ram_mem2_255_16,
         p_wishbone_bd_ram_mem2_255_17, p_wishbone_bd_ram_mem2_255_18,
         p_wishbone_bd_ram_mem2_255_19, p_wishbone_bd_ram_mem2_255_20,
         p_wishbone_bd_ram_mem2_255_21, p_wishbone_bd_ram_mem2_255_22,
         p_wishbone_bd_ram_mem2_255_23, p_wishbone_bd_ram_mem3_0_24,
         p_wishbone_bd_ram_mem3_0_25, p_wishbone_bd_ram_mem3_0_26,
         p_wishbone_bd_ram_mem3_0_27, p_wishbone_bd_ram_mem3_0_28,
         p_wishbone_bd_ram_mem3_0_29, p_wishbone_bd_ram_mem3_0_30,
         p_wishbone_bd_ram_mem3_0_31, p_wishbone_bd_ram_mem3_1_24,
         p_wishbone_bd_ram_mem3_1_25, p_wishbone_bd_ram_mem3_1_26,
         p_wishbone_bd_ram_mem3_1_27, p_wishbone_bd_ram_mem3_1_28,
         p_wishbone_bd_ram_mem3_1_29, p_wishbone_bd_ram_mem3_1_30,
         p_wishbone_bd_ram_mem3_1_31, p_wishbone_bd_ram_mem3_2_24,
         p_wishbone_bd_ram_mem3_2_25, p_wishbone_bd_ram_mem3_2_26,
         p_wishbone_bd_ram_mem3_2_27, p_wishbone_bd_ram_mem3_2_28,
         p_wishbone_bd_ram_mem3_2_29, p_wishbone_bd_ram_mem3_2_30,
         p_wishbone_bd_ram_mem3_2_31, p_wishbone_bd_ram_mem3_3_24,
         p_wishbone_bd_ram_mem3_3_25, p_wishbone_bd_ram_mem3_3_26,
         p_wishbone_bd_ram_mem3_3_27, p_wishbone_bd_ram_mem3_3_28,
         p_wishbone_bd_ram_mem3_3_29, p_wishbone_bd_ram_mem3_3_30,
         p_wishbone_bd_ram_mem3_3_31, p_wishbone_bd_ram_mem3_4_24,
         p_wishbone_bd_ram_mem3_4_25, p_wishbone_bd_ram_mem3_4_26,
         p_wishbone_bd_ram_mem3_4_27, p_wishbone_bd_ram_mem3_4_28,
         p_wishbone_bd_ram_mem3_4_29, p_wishbone_bd_ram_mem3_4_30,
         p_wishbone_bd_ram_mem3_4_31, p_wishbone_bd_ram_mem3_5_24,
         p_wishbone_bd_ram_mem3_5_25, p_wishbone_bd_ram_mem3_5_26,
         p_wishbone_bd_ram_mem3_5_27, p_wishbone_bd_ram_mem3_5_28,
         p_wishbone_bd_ram_mem3_5_29, p_wishbone_bd_ram_mem3_5_30,
         p_wishbone_bd_ram_mem3_5_31, p_wishbone_bd_ram_mem3_6_24,
         p_wishbone_bd_ram_mem3_6_25, p_wishbone_bd_ram_mem3_6_26,
         p_wishbone_bd_ram_mem3_6_27, p_wishbone_bd_ram_mem3_6_28,
         p_wishbone_bd_ram_mem3_6_29, p_wishbone_bd_ram_mem3_6_30,
         p_wishbone_bd_ram_mem3_6_31, p_wishbone_bd_ram_mem3_7_24,
         p_wishbone_bd_ram_mem3_7_25, p_wishbone_bd_ram_mem3_7_26,
         p_wishbone_bd_ram_mem3_7_27, p_wishbone_bd_ram_mem3_7_28,
         p_wishbone_bd_ram_mem3_7_29, p_wishbone_bd_ram_mem3_7_30,
         p_wishbone_bd_ram_mem3_7_31, p_wishbone_bd_ram_mem3_8_24,
         p_wishbone_bd_ram_mem3_8_25, p_wishbone_bd_ram_mem3_8_26,
         p_wishbone_bd_ram_mem3_8_27, p_wishbone_bd_ram_mem3_8_28,
         p_wishbone_bd_ram_mem3_8_29, p_wishbone_bd_ram_mem3_8_30,
         p_wishbone_bd_ram_mem3_8_31, p_wishbone_bd_ram_mem3_9_24,
         p_wishbone_bd_ram_mem3_9_25, p_wishbone_bd_ram_mem3_9_26,
         p_wishbone_bd_ram_mem3_9_27, p_wishbone_bd_ram_mem3_9_28,
         p_wishbone_bd_ram_mem3_9_29, p_wishbone_bd_ram_mem3_9_30,
         p_wishbone_bd_ram_mem3_9_31, p_wishbone_bd_ram_mem3_10_24,
         p_wishbone_bd_ram_mem3_10_25, p_wishbone_bd_ram_mem3_10_26,
         p_wishbone_bd_ram_mem3_10_27, p_wishbone_bd_ram_mem3_10_28,
         p_wishbone_bd_ram_mem3_10_29, p_wishbone_bd_ram_mem3_10_30,
         p_wishbone_bd_ram_mem3_10_31, p_wishbone_bd_ram_mem3_11_24,
         p_wishbone_bd_ram_mem3_11_25, p_wishbone_bd_ram_mem3_11_26,
         p_wishbone_bd_ram_mem3_11_27, p_wishbone_bd_ram_mem3_11_28,
         p_wishbone_bd_ram_mem3_11_29, p_wishbone_bd_ram_mem3_11_30,
         p_wishbone_bd_ram_mem3_11_31, p_wishbone_bd_ram_mem3_12_24,
         p_wishbone_bd_ram_mem3_12_25, p_wishbone_bd_ram_mem3_12_26,
         p_wishbone_bd_ram_mem3_12_27, p_wishbone_bd_ram_mem3_12_28,
         p_wishbone_bd_ram_mem3_12_29, p_wishbone_bd_ram_mem3_12_30,
         p_wishbone_bd_ram_mem3_12_31, p_wishbone_bd_ram_mem3_13_24,
         p_wishbone_bd_ram_mem3_13_25, p_wishbone_bd_ram_mem3_13_26,
         p_wishbone_bd_ram_mem3_13_27, p_wishbone_bd_ram_mem3_13_28,
         p_wishbone_bd_ram_mem3_13_29, p_wishbone_bd_ram_mem3_13_30,
         p_wishbone_bd_ram_mem3_13_31, p_wishbone_bd_ram_mem3_14_24,
         p_wishbone_bd_ram_mem3_14_25, p_wishbone_bd_ram_mem3_14_26,
         p_wishbone_bd_ram_mem3_14_27, p_wishbone_bd_ram_mem3_14_28,
         p_wishbone_bd_ram_mem3_14_29, p_wishbone_bd_ram_mem3_14_30,
         p_wishbone_bd_ram_mem3_14_31, p_wishbone_bd_ram_mem3_15_24,
         p_wishbone_bd_ram_mem3_15_25, p_wishbone_bd_ram_mem3_15_26,
         p_wishbone_bd_ram_mem3_15_27, p_wishbone_bd_ram_mem3_15_28,
         p_wishbone_bd_ram_mem3_15_29, p_wishbone_bd_ram_mem3_15_30,
         p_wishbone_bd_ram_mem3_15_31, p_wishbone_bd_ram_mem3_16_24,
         p_wishbone_bd_ram_mem3_16_25, p_wishbone_bd_ram_mem3_16_26,
         p_wishbone_bd_ram_mem3_16_27, p_wishbone_bd_ram_mem3_16_28,
         p_wishbone_bd_ram_mem3_16_29, p_wishbone_bd_ram_mem3_16_30,
         p_wishbone_bd_ram_mem3_16_31, p_wishbone_bd_ram_mem3_17_24,
         p_wishbone_bd_ram_mem3_17_25, p_wishbone_bd_ram_mem3_17_26,
         p_wishbone_bd_ram_mem3_17_27, p_wishbone_bd_ram_mem3_17_28,
         p_wishbone_bd_ram_mem3_17_29, p_wishbone_bd_ram_mem3_17_30,
         p_wishbone_bd_ram_mem3_17_31, p_wishbone_bd_ram_mem3_18_24,
         p_wishbone_bd_ram_mem3_18_25, p_wishbone_bd_ram_mem3_18_26,
         p_wishbone_bd_ram_mem3_18_27, p_wishbone_bd_ram_mem3_18_28,
         p_wishbone_bd_ram_mem3_18_29, p_wishbone_bd_ram_mem3_18_30,
         p_wishbone_bd_ram_mem3_18_31, p_wishbone_bd_ram_mem3_19_24,
         p_wishbone_bd_ram_mem3_19_25, p_wishbone_bd_ram_mem3_19_26,
         p_wishbone_bd_ram_mem3_19_27, p_wishbone_bd_ram_mem3_19_28,
         p_wishbone_bd_ram_mem3_19_29, p_wishbone_bd_ram_mem3_19_30,
         p_wishbone_bd_ram_mem3_19_31, p_wishbone_bd_ram_mem3_20_24,
         p_wishbone_bd_ram_mem3_20_25, p_wishbone_bd_ram_mem3_20_26,
         p_wishbone_bd_ram_mem3_20_27, p_wishbone_bd_ram_mem3_20_28,
         p_wishbone_bd_ram_mem3_20_29, p_wishbone_bd_ram_mem3_20_30,
         p_wishbone_bd_ram_mem3_20_31, p_wishbone_bd_ram_mem3_21_24,
         p_wishbone_bd_ram_mem3_21_25, p_wishbone_bd_ram_mem3_21_26,
         p_wishbone_bd_ram_mem3_21_27, p_wishbone_bd_ram_mem3_21_28,
         p_wishbone_bd_ram_mem3_21_29, p_wishbone_bd_ram_mem3_21_30,
         p_wishbone_bd_ram_mem3_21_31, p_wishbone_bd_ram_mem3_22_24,
         p_wishbone_bd_ram_mem3_22_25, p_wishbone_bd_ram_mem3_22_26,
         p_wishbone_bd_ram_mem3_22_27, p_wishbone_bd_ram_mem3_22_28,
         p_wishbone_bd_ram_mem3_22_29, p_wishbone_bd_ram_mem3_22_30,
         p_wishbone_bd_ram_mem3_22_31, p_wishbone_bd_ram_mem3_23_24,
         p_wishbone_bd_ram_mem3_23_25, p_wishbone_bd_ram_mem3_23_26,
         p_wishbone_bd_ram_mem3_23_27, p_wishbone_bd_ram_mem3_23_28,
         p_wishbone_bd_ram_mem3_23_29, p_wishbone_bd_ram_mem3_23_30,
         p_wishbone_bd_ram_mem3_23_31, p_wishbone_bd_ram_mem3_24_24,
         p_wishbone_bd_ram_mem3_24_25, p_wishbone_bd_ram_mem3_24_26,
         p_wishbone_bd_ram_mem3_24_27, p_wishbone_bd_ram_mem3_24_28,
         p_wishbone_bd_ram_mem3_24_29, p_wishbone_bd_ram_mem3_24_30,
         p_wishbone_bd_ram_mem3_24_31, p_wishbone_bd_ram_mem3_25_24,
         p_wishbone_bd_ram_mem3_25_25, p_wishbone_bd_ram_mem3_25_26,
         p_wishbone_bd_ram_mem3_25_27, p_wishbone_bd_ram_mem3_25_28,
         p_wishbone_bd_ram_mem3_25_29, p_wishbone_bd_ram_mem3_25_30,
         p_wishbone_bd_ram_mem3_25_31, p_wishbone_bd_ram_mem3_26_24,
         p_wishbone_bd_ram_mem3_26_25, p_wishbone_bd_ram_mem3_26_26,
         p_wishbone_bd_ram_mem3_26_27, p_wishbone_bd_ram_mem3_26_28,
         p_wishbone_bd_ram_mem3_26_29, p_wishbone_bd_ram_mem3_26_30,
         p_wishbone_bd_ram_mem3_26_31, p_wishbone_bd_ram_mem3_27_24,
         p_wishbone_bd_ram_mem3_27_25, p_wishbone_bd_ram_mem3_27_26,
         p_wishbone_bd_ram_mem3_27_27, p_wishbone_bd_ram_mem3_27_28,
         p_wishbone_bd_ram_mem3_27_29, p_wishbone_bd_ram_mem3_27_30,
         p_wishbone_bd_ram_mem3_27_31, p_wishbone_bd_ram_mem3_28_24,
         p_wishbone_bd_ram_mem3_28_25, p_wishbone_bd_ram_mem3_28_26,
         p_wishbone_bd_ram_mem3_28_27, p_wishbone_bd_ram_mem3_28_28,
         p_wishbone_bd_ram_mem3_28_29, p_wishbone_bd_ram_mem3_28_30,
         p_wishbone_bd_ram_mem3_28_31, p_wishbone_bd_ram_mem3_29_24,
         p_wishbone_bd_ram_mem3_29_25, p_wishbone_bd_ram_mem3_29_26,
         p_wishbone_bd_ram_mem3_29_27, p_wishbone_bd_ram_mem3_29_28,
         p_wishbone_bd_ram_mem3_29_29, p_wishbone_bd_ram_mem3_29_30,
         p_wishbone_bd_ram_mem3_29_31, p_wishbone_bd_ram_mem3_30_24,
         p_wishbone_bd_ram_mem3_30_25, p_wishbone_bd_ram_mem3_30_26,
         p_wishbone_bd_ram_mem3_30_27, p_wishbone_bd_ram_mem3_30_28,
         p_wishbone_bd_ram_mem3_30_29, p_wishbone_bd_ram_mem3_30_30,
         p_wishbone_bd_ram_mem3_30_31, p_wishbone_bd_ram_mem3_31_24,
         p_wishbone_bd_ram_mem3_31_25, p_wishbone_bd_ram_mem3_31_26,
         p_wishbone_bd_ram_mem3_31_27, p_wishbone_bd_ram_mem3_31_28,
         p_wishbone_bd_ram_mem3_31_29, p_wishbone_bd_ram_mem3_31_30,
         p_wishbone_bd_ram_mem3_31_31, p_wishbone_bd_ram_mem3_32_24,
         p_wishbone_bd_ram_mem3_32_25, p_wishbone_bd_ram_mem3_32_26,
         p_wishbone_bd_ram_mem3_32_27, p_wishbone_bd_ram_mem3_32_28,
         p_wishbone_bd_ram_mem3_32_29, p_wishbone_bd_ram_mem3_32_30,
         p_wishbone_bd_ram_mem3_32_31, p_wishbone_bd_ram_mem3_33_24,
         p_wishbone_bd_ram_mem3_33_25, p_wishbone_bd_ram_mem3_33_26,
         p_wishbone_bd_ram_mem3_33_27, p_wishbone_bd_ram_mem3_33_28,
         p_wishbone_bd_ram_mem3_33_29, p_wishbone_bd_ram_mem3_33_30,
         p_wishbone_bd_ram_mem3_33_31, p_wishbone_bd_ram_mem3_34_24,
         p_wishbone_bd_ram_mem3_34_25, p_wishbone_bd_ram_mem3_34_26,
         p_wishbone_bd_ram_mem3_34_27, p_wishbone_bd_ram_mem3_34_28,
         p_wishbone_bd_ram_mem3_34_29, p_wishbone_bd_ram_mem3_34_30,
         p_wishbone_bd_ram_mem3_34_31, p_wishbone_bd_ram_mem3_35_24,
         p_wishbone_bd_ram_mem3_35_25, p_wishbone_bd_ram_mem3_35_26,
         p_wishbone_bd_ram_mem3_35_27, p_wishbone_bd_ram_mem3_35_28,
         p_wishbone_bd_ram_mem3_35_29, p_wishbone_bd_ram_mem3_35_30,
         p_wishbone_bd_ram_mem3_35_31, p_wishbone_bd_ram_mem3_36_24,
         p_wishbone_bd_ram_mem3_36_25, p_wishbone_bd_ram_mem3_36_26,
         p_wishbone_bd_ram_mem3_36_27, p_wishbone_bd_ram_mem3_36_28,
         p_wishbone_bd_ram_mem3_36_29, p_wishbone_bd_ram_mem3_36_30,
         p_wishbone_bd_ram_mem3_36_31, p_wishbone_bd_ram_mem3_37_24,
         p_wishbone_bd_ram_mem3_37_25, p_wishbone_bd_ram_mem3_37_26,
         p_wishbone_bd_ram_mem3_37_27, p_wishbone_bd_ram_mem3_37_28,
         p_wishbone_bd_ram_mem3_37_29, p_wishbone_bd_ram_mem3_37_30,
         p_wishbone_bd_ram_mem3_37_31, p_wishbone_bd_ram_mem3_38_24,
         p_wishbone_bd_ram_mem3_38_25, p_wishbone_bd_ram_mem3_38_26,
         p_wishbone_bd_ram_mem3_38_27, p_wishbone_bd_ram_mem3_38_28,
         p_wishbone_bd_ram_mem3_38_29, p_wishbone_bd_ram_mem3_38_30,
         p_wishbone_bd_ram_mem3_38_31, p_wishbone_bd_ram_mem3_39_24,
         p_wishbone_bd_ram_mem3_39_25, p_wishbone_bd_ram_mem3_39_26,
         p_wishbone_bd_ram_mem3_39_27, p_wishbone_bd_ram_mem3_39_28,
         p_wishbone_bd_ram_mem3_39_29, p_wishbone_bd_ram_mem3_39_30,
         p_wishbone_bd_ram_mem3_39_31, p_wishbone_bd_ram_mem3_40_24,
         p_wishbone_bd_ram_mem3_40_25, p_wishbone_bd_ram_mem3_40_26,
         p_wishbone_bd_ram_mem3_40_27, p_wishbone_bd_ram_mem3_40_28,
         p_wishbone_bd_ram_mem3_40_29, p_wishbone_bd_ram_mem3_40_30,
         p_wishbone_bd_ram_mem3_40_31, p_wishbone_bd_ram_mem3_41_24,
         p_wishbone_bd_ram_mem3_41_25, p_wishbone_bd_ram_mem3_41_26,
         p_wishbone_bd_ram_mem3_41_27, p_wishbone_bd_ram_mem3_41_28,
         p_wishbone_bd_ram_mem3_41_29, p_wishbone_bd_ram_mem3_41_30,
         p_wishbone_bd_ram_mem3_41_31, p_wishbone_bd_ram_mem3_42_24,
         p_wishbone_bd_ram_mem3_42_25, p_wishbone_bd_ram_mem3_42_26,
         p_wishbone_bd_ram_mem3_42_27, p_wishbone_bd_ram_mem3_42_28,
         p_wishbone_bd_ram_mem3_42_29, p_wishbone_bd_ram_mem3_42_30,
         p_wishbone_bd_ram_mem3_42_31, p_wishbone_bd_ram_mem3_43_24,
         p_wishbone_bd_ram_mem3_43_25, p_wishbone_bd_ram_mem3_43_26,
         p_wishbone_bd_ram_mem3_43_27, p_wishbone_bd_ram_mem3_43_28,
         p_wishbone_bd_ram_mem3_43_29, p_wishbone_bd_ram_mem3_43_30,
         p_wishbone_bd_ram_mem3_43_31, p_wishbone_bd_ram_mem3_44_24,
         p_wishbone_bd_ram_mem3_44_25, p_wishbone_bd_ram_mem3_44_26,
         p_wishbone_bd_ram_mem3_44_27, p_wishbone_bd_ram_mem3_44_28,
         p_wishbone_bd_ram_mem3_44_29, p_wishbone_bd_ram_mem3_44_30,
         p_wishbone_bd_ram_mem3_44_31, p_wishbone_bd_ram_mem3_45_24,
         p_wishbone_bd_ram_mem3_45_25, p_wishbone_bd_ram_mem3_45_26,
         p_wishbone_bd_ram_mem3_45_27, p_wishbone_bd_ram_mem3_45_28,
         p_wishbone_bd_ram_mem3_45_29, p_wishbone_bd_ram_mem3_45_30,
         p_wishbone_bd_ram_mem3_45_31, p_wishbone_bd_ram_mem3_46_24,
         p_wishbone_bd_ram_mem3_46_25, p_wishbone_bd_ram_mem3_46_26,
         p_wishbone_bd_ram_mem3_46_27, p_wishbone_bd_ram_mem3_46_28,
         p_wishbone_bd_ram_mem3_46_29, p_wishbone_bd_ram_mem3_46_30,
         p_wishbone_bd_ram_mem3_46_31, p_wishbone_bd_ram_mem3_47_24,
         p_wishbone_bd_ram_mem3_47_25, p_wishbone_bd_ram_mem3_47_26,
         p_wishbone_bd_ram_mem3_47_27, p_wishbone_bd_ram_mem3_47_28,
         p_wishbone_bd_ram_mem3_47_29, p_wishbone_bd_ram_mem3_47_30,
         p_wishbone_bd_ram_mem3_47_31, p_wishbone_bd_ram_mem3_48_24,
         p_wishbone_bd_ram_mem3_48_25, p_wishbone_bd_ram_mem3_48_26,
         p_wishbone_bd_ram_mem3_48_27, p_wishbone_bd_ram_mem3_48_28,
         p_wishbone_bd_ram_mem3_48_29, p_wishbone_bd_ram_mem3_48_30,
         p_wishbone_bd_ram_mem3_48_31, p_wishbone_bd_ram_mem3_49_24,
         p_wishbone_bd_ram_mem3_49_25, p_wishbone_bd_ram_mem3_49_26,
         p_wishbone_bd_ram_mem3_49_27, p_wishbone_bd_ram_mem3_49_28,
         p_wishbone_bd_ram_mem3_49_29, p_wishbone_bd_ram_mem3_49_30,
         p_wishbone_bd_ram_mem3_49_31, p_wishbone_bd_ram_mem3_50_24,
         p_wishbone_bd_ram_mem3_50_25, p_wishbone_bd_ram_mem3_50_26,
         p_wishbone_bd_ram_mem3_50_27, p_wishbone_bd_ram_mem3_50_28,
         p_wishbone_bd_ram_mem3_50_29, p_wishbone_bd_ram_mem3_50_30,
         p_wishbone_bd_ram_mem3_50_31, p_wishbone_bd_ram_mem3_51_24,
         p_wishbone_bd_ram_mem3_51_25, p_wishbone_bd_ram_mem3_51_26,
         p_wishbone_bd_ram_mem3_51_27, p_wishbone_bd_ram_mem3_51_28,
         p_wishbone_bd_ram_mem3_51_29, p_wishbone_bd_ram_mem3_51_30,
         p_wishbone_bd_ram_mem3_51_31, p_wishbone_bd_ram_mem3_52_24,
         p_wishbone_bd_ram_mem3_52_25, p_wishbone_bd_ram_mem3_52_26,
         p_wishbone_bd_ram_mem3_52_27, p_wishbone_bd_ram_mem3_52_28,
         p_wishbone_bd_ram_mem3_52_29, p_wishbone_bd_ram_mem3_52_30,
         p_wishbone_bd_ram_mem3_52_31, p_wishbone_bd_ram_mem3_53_24,
         p_wishbone_bd_ram_mem3_53_25, p_wishbone_bd_ram_mem3_53_26,
         p_wishbone_bd_ram_mem3_53_27, p_wishbone_bd_ram_mem3_53_28,
         p_wishbone_bd_ram_mem3_53_29, p_wishbone_bd_ram_mem3_53_30,
         p_wishbone_bd_ram_mem3_53_31, p_wishbone_bd_ram_mem3_54_24,
         p_wishbone_bd_ram_mem3_54_25, p_wishbone_bd_ram_mem3_54_26,
         p_wishbone_bd_ram_mem3_54_27, p_wishbone_bd_ram_mem3_54_28,
         p_wishbone_bd_ram_mem3_54_29, p_wishbone_bd_ram_mem3_54_30,
         p_wishbone_bd_ram_mem3_54_31, p_wishbone_bd_ram_mem3_55_24,
         p_wishbone_bd_ram_mem3_55_25, p_wishbone_bd_ram_mem3_55_26,
         p_wishbone_bd_ram_mem3_55_27, p_wishbone_bd_ram_mem3_55_28,
         p_wishbone_bd_ram_mem3_55_29, p_wishbone_bd_ram_mem3_55_30,
         p_wishbone_bd_ram_mem3_55_31, p_wishbone_bd_ram_mem3_56_24,
         p_wishbone_bd_ram_mem3_56_25, p_wishbone_bd_ram_mem3_56_26,
         p_wishbone_bd_ram_mem3_56_27, p_wishbone_bd_ram_mem3_56_28,
         p_wishbone_bd_ram_mem3_56_29, p_wishbone_bd_ram_mem3_56_30,
         p_wishbone_bd_ram_mem3_56_31, p_wishbone_bd_ram_mem3_57_24,
         p_wishbone_bd_ram_mem3_57_25, p_wishbone_bd_ram_mem3_57_26,
         p_wishbone_bd_ram_mem3_57_27, p_wishbone_bd_ram_mem3_57_28,
         p_wishbone_bd_ram_mem3_57_29, p_wishbone_bd_ram_mem3_57_30,
         p_wishbone_bd_ram_mem3_57_31, p_wishbone_bd_ram_mem3_58_24,
         p_wishbone_bd_ram_mem3_58_25, p_wishbone_bd_ram_mem3_58_26,
         p_wishbone_bd_ram_mem3_58_27, p_wishbone_bd_ram_mem3_58_28,
         p_wishbone_bd_ram_mem3_58_29, p_wishbone_bd_ram_mem3_58_30,
         p_wishbone_bd_ram_mem3_58_31, p_wishbone_bd_ram_mem3_59_24,
         p_wishbone_bd_ram_mem3_59_25, p_wishbone_bd_ram_mem3_59_26,
         p_wishbone_bd_ram_mem3_59_27, p_wishbone_bd_ram_mem3_59_28,
         p_wishbone_bd_ram_mem3_59_29, p_wishbone_bd_ram_mem3_59_30,
         p_wishbone_bd_ram_mem3_59_31, p_wishbone_bd_ram_mem3_60_24,
         p_wishbone_bd_ram_mem3_60_25, p_wishbone_bd_ram_mem3_60_26,
         p_wishbone_bd_ram_mem3_60_27, p_wishbone_bd_ram_mem3_60_28,
         p_wishbone_bd_ram_mem3_60_29, p_wishbone_bd_ram_mem3_60_30,
         p_wishbone_bd_ram_mem3_60_31, p_wishbone_bd_ram_mem3_61_24,
         p_wishbone_bd_ram_mem3_61_25, p_wishbone_bd_ram_mem3_61_26,
         p_wishbone_bd_ram_mem3_61_27, p_wishbone_bd_ram_mem3_61_28,
         p_wishbone_bd_ram_mem3_61_29, p_wishbone_bd_ram_mem3_61_30,
         p_wishbone_bd_ram_mem3_61_31, p_wishbone_bd_ram_mem3_62_24,
         p_wishbone_bd_ram_mem3_62_25, p_wishbone_bd_ram_mem3_62_26,
         p_wishbone_bd_ram_mem3_62_27, p_wishbone_bd_ram_mem3_62_28,
         p_wishbone_bd_ram_mem3_62_29, p_wishbone_bd_ram_mem3_62_30,
         p_wishbone_bd_ram_mem3_62_31, p_wishbone_bd_ram_mem3_63_24,
         p_wishbone_bd_ram_mem3_63_25, p_wishbone_bd_ram_mem3_63_26,
         p_wishbone_bd_ram_mem3_63_27, p_wishbone_bd_ram_mem3_63_28,
         p_wishbone_bd_ram_mem3_63_29, p_wishbone_bd_ram_mem3_63_30,
         p_wishbone_bd_ram_mem3_63_31, p_wishbone_bd_ram_mem3_64_24,
         p_wishbone_bd_ram_mem3_64_25, p_wishbone_bd_ram_mem3_64_26,
         p_wishbone_bd_ram_mem3_64_27, p_wishbone_bd_ram_mem3_64_28,
         p_wishbone_bd_ram_mem3_64_29, p_wishbone_bd_ram_mem3_64_30,
         p_wishbone_bd_ram_mem3_64_31, p_wishbone_bd_ram_mem3_65_24,
         p_wishbone_bd_ram_mem3_65_25, p_wishbone_bd_ram_mem3_65_26,
         p_wishbone_bd_ram_mem3_65_27, p_wishbone_bd_ram_mem3_65_28,
         p_wishbone_bd_ram_mem3_65_29, p_wishbone_bd_ram_mem3_65_30,
         p_wishbone_bd_ram_mem3_65_31, p_wishbone_bd_ram_mem3_66_24,
         p_wishbone_bd_ram_mem3_66_25, p_wishbone_bd_ram_mem3_66_26,
         p_wishbone_bd_ram_mem3_66_27, p_wishbone_bd_ram_mem3_66_28,
         p_wishbone_bd_ram_mem3_66_29, p_wishbone_bd_ram_mem3_66_30,
         p_wishbone_bd_ram_mem3_66_31, p_wishbone_bd_ram_mem3_67_24,
         p_wishbone_bd_ram_mem3_67_25, p_wishbone_bd_ram_mem3_67_26,
         p_wishbone_bd_ram_mem3_67_27, p_wishbone_bd_ram_mem3_67_28,
         p_wishbone_bd_ram_mem3_67_29, p_wishbone_bd_ram_mem3_67_30,
         p_wishbone_bd_ram_mem3_67_31, p_wishbone_bd_ram_mem3_68_24,
         p_wishbone_bd_ram_mem3_68_25, p_wishbone_bd_ram_mem3_68_26,
         p_wishbone_bd_ram_mem3_68_27, p_wishbone_bd_ram_mem3_68_28,
         p_wishbone_bd_ram_mem3_68_29, p_wishbone_bd_ram_mem3_68_30,
         p_wishbone_bd_ram_mem3_68_31, p_wishbone_bd_ram_mem3_69_24,
         p_wishbone_bd_ram_mem3_69_25, p_wishbone_bd_ram_mem3_69_26,
         p_wishbone_bd_ram_mem3_69_27, p_wishbone_bd_ram_mem3_69_28,
         p_wishbone_bd_ram_mem3_69_29, p_wishbone_bd_ram_mem3_69_30,
         p_wishbone_bd_ram_mem3_69_31, p_wishbone_bd_ram_mem3_70_24,
         p_wishbone_bd_ram_mem3_70_25, p_wishbone_bd_ram_mem3_70_26,
         p_wishbone_bd_ram_mem3_70_27, p_wishbone_bd_ram_mem3_70_28,
         p_wishbone_bd_ram_mem3_70_29, p_wishbone_bd_ram_mem3_70_30,
         p_wishbone_bd_ram_mem3_70_31, p_wishbone_bd_ram_mem3_71_24,
         p_wishbone_bd_ram_mem3_71_25, p_wishbone_bd_ram_mem3_71_26,
         p_wishbone_bd_ram_mem3_71_27, p_wishbone_bd_ram_mem3_71_28,
         p_wishbone_bd_ram_mem3_71_29, p_wishbone_bd_ram_mem3_71_30,
         p_wishbone_bd_ram_mem3_71_31, p_wishbone_bd_ram_mem3_72_24,
         p_wishbone_bd_ram_mem3_72_25, p_wishbone_bd_ram_mem3_72_26,
         p_wishbone_bd_ram_mem3_72_27, p_wishbone_bd_ram_mem3_72_28,
         p_wishbone_bd_ram_mem3_72_29, p_wishbone_bd_ram_mem3_72_30,
         p_wishbone_bd_ram_mem3_72_31, p_wishbone_bd_ram_mem3_73_24,
         p_wishbone_bd_ram_mem3_73_25, p_wishbone_bd_ram_mem3_73_26,
         p_wishbone_bd_ram_mem3_73_27, p_wishbone_bd_ram_mem3_73_28,
         p_wishbone_bd_ram_mem3_73_29, p_wishbone_bd_ram_mem3_73_30,
         p_wishbone_bd_ram_mem3_73_31, p_wishbone_bd_ram_mem3_74_24,
         p_wishbone_bd_ram_mem3_74_25, p_wishbone_bd_ram_mem3_74_26,
         p_wishbone_bd_ram_mem3_74_27, p_wishbone_bd_ram_mem3_74_28,
         p_wishbone_bd_ram_mem3_74_29, p_wishbone_bd_ram_mem3_74_30,
         p_wishbone_bd_ram_mem3_74_31, p_wishbone_bd_ram_mem3_75_24,
         p_wishbone_bd_ram_mem3_75_25, p_wishbone_bd_ram_mem3_75_26,
         p_wishbone_bd_ram_mem3_75_27, p_wishbone_bd_ram_mem3_75_28,
         p_wishbone_bd_ram_mem3_75_29, p_wishbone_bd_ram_mem3_75_30,
         p_wishbone_bd_ram_mem3_75_31, p_wishbone_bd_ram_mem3_76_24,
         p_wishbone_bd_ram_mem3_76_25, p_wishbone_bd_ram_mem3_76_26,
         p_wishbone_bd_ram_mem3_76_27, p_wishbone_bd_ram_mem3_76_28,
         p_wishbone_bd_ram_mem3_76_29, p_wishbone_bd_ram_mem3_76_30,
         p_wishbone_bd_ram_mem3_76_31, p_wishbone_bd_ram_mem3_77_24,
         p_wishbone_bd_ram_mem3_77_25, p_wishbone_bd_ram_mem3_77_26,
         p_wishbone_bd_ram_mem3_77_27, p_wishbone_bd_ram_mem3_77_28,
         p_wishbone_bd_ram_mem3_77_29, p_wishbone_bd_ram_mem3_77_30,
         p_wishbone_bd_ram_mem3_77_31, p_wishbone_bd_ram_mem3_78_24,
         p_wishbone_bd_ram_mem3_78_25, p_wishbone_bd_ram_mem3_78_26,
         p_wishbone_bd_ram_mem3_78_27, p_wishbone_bd_ram_mem3_78_28,
         p_wishbone_bd_ram_mem3_78_29, p_wishbone_bd_ram_mem3_78_30,
         p_wishbone_bd_ram_mem3_78_31, p_wishbone_bd_ram_mem3_79_24,
         p_wishbone_bd_ram_mem3_79_25, p_wishbone_bd_ram_mem3_79_26,
         p_wishbone_bd_ram_mem3_79_27, p_wishbone_bd_ram_mem3_79_28,
         p_wishbone_bd_ram_mem3_79_29, p_wishbone_bd_ram_mem3_79_30,
         p_wishbone_bd_ram_mem3_79_31, p_wishbone_bd_ram_mem3_80_24,
         p_wishbone_bd_ram_mem3_80_25, p_wishbone_bd_ram_mem3_80_26,
         p_wishbone_bd_ram_mem3_80_27, p_wishbone_bd_ram_mem3_80_28,
         p_wishbone_bd_ram_mem3_80_29, p_wishbone_bd_ram_mem3_80_30,
         p_wishbone_bd_ram_mem3_80_31, p_wishbone_bd_ram_mem3_81_24,
         p_wishbone_bd_ram_mem3_81_25, p_wishbone_bd_ram_mem3_81_26,
         p_wishbone_bd_ram_mem3_81_27, p_wishbone_bd_ram_mem3_81_28,
         p_wishbone_bd_ram_mem3_81_29, p_wishbone_bd_ram_mem3_81_30,
         p_wishbone_bd_ram_mem3_81_31, p_wishbone_bd_ram_mem3_82_24,
         p_wishbone_bd_ram_mem3_82_25, p_wishbone_bd_ram_mem3_82_26,
         p_wishbone_bd_ram_mem3_82_27, p_wishbone_bd_ram_mem3_82_28,
         p_wishbone_bd_ram_mem3_82_29, p_wishbone_bd_ram_mem3_82_30,
         p_wishbone_bd_ram_mem3_82_31, p_wishbone_bd_ram_mem3_83_24,
         p_wishbone_bd_ram_mem3_83_25, p_wishbone_bd_ram_mem3_83_26,
         p_wishbone_bd_ram_mem3_83_27, p_wishbone_bd_ram_mem3_83_28,
         p_wishbone_bd_ram_mem3_83_29, p_wishbone_bd_ram_mem3_83_30,
         p_wishbone_bd_ram_mem3_83_31, p_wishbone_bd_ram_mem3_84_24,
         p_wishbone_bd_ram_mem3_84_25, p_wishbone_bd_ram_mem3_84_26,
         p_wishbone_bd_ram_mem3_84_27, p_wishbone_bd_ram_mem3_84_28,
         p_wishbone_bd_ram_mem3_84_29, p_wishbone_bd_ram_mem3_84_30,
         p_wishbone_bd_ram_mem3_84_31, p_wishbone_bd_ram_mem3_85_24,
         p_wishbone_bd_ram_mem3_85_25, p_wishbone_bd_ram_mem3_85_26,
         p_wishbone_bd_ram_mem3_85_27, p_wishbone_bd_ram_mem3_85_28,
         p_wishbone_bd_ram_mem3_85_29, p_wishbone_bd_ram_mem3_85_30,
         p_wishbone_bd_ram_mem3_85_31, p_wishbone_bd_ram_mem3_86_24,
         p_wishbone_bd_ram_mem3_86_25, p_wishbone_bd_ram_mem3_86_26,
         p_wishbone_bd_ram_mem3_86_27, p_wishbone_bd_ram_mem3_86_28,
         p_wishbone_bd_ram_mem3_86_29, p_wishbone_bd_ram_mem3_86_30,
         p_wishbone_bd_ram_mem3_86_31, p_wishbone_bd_ram_mem3_87_24,
         p_wishbone_bd_ram_mem3_87_25, p_wishbone_bd_ram_mem3_87_26,
         p_wishbone_bd_ram_mem3_87_27, p_wishbone_bd_ram_mem3_87_28,
         p_wishbone_bd_ram_mem3_87_29, p_wishbone_bd_ram_mem3_87_30,
         p_wishbone_bd_ram_mem3_87_31, p_wishbone_bd_ram_mem3_88_24,
         p_wishbone_bd_ram_mem3_88_25, p_wishbone_bd_ram_mem3_88_26,
         p_wishbone_bd_ram_mem3_88_27, p_wishbone_bd_ram_mem3_88_28,
         p_wishbone_bd_ram_mem3_88_29, p_wishbone_bd_ram_mem3_88_30,
         p_wishbone_bd_ram_mem3_88_31, p_wishbone_bd_ram_mem3_89_24,
         p_wishbone_bd_ram_mem3_89_25, p_wishbone_bd_ram_mem3_89_26,
         p_wishbone_bd_ram_mem3_89_27, p_wishbone_bd_ram_mem3_89_28,
         p_wishbone_bd_ram_mem3_89_29, p_wishbone_bd_ram_mem3_89_30,
         p_wishbone_bd_ram_mem3_89_31, p_wishbone_bd_ram_mem3_90_24,
         p_wishbone_bd_ram_mem3_90_25, p_wishbone_bd_ram_mem3_90_26,
         p_wishbone_bd_ram_mem3_90_27, p_wishbone_bd_ram_mem3_90_28,
         p_wishbone_bd_ram_mem3_90_29, p_wishbone_bd_ram_mem3_90_30,
         p_wishbone_bd_ram_mem3_90_31, p_wishbone_bd_ram_mem3_91_24,
         p_wishbone_bd_ram_mem3_91_25, p_wishbone_bd_ram_mem3_91_26,
         p_wishbone_bd_ram_mem3_91_27, p_wishbone_bd_ram_mem3_91_28,
         p_wishbone_bd_ram_mem3_91_29, p_wishbone_bd_ram_mem3_91_30,
         p_wishbone_bd_ram_mem3_91_31, p_wishbone_bd_ram_mem3_92_24,
         p_wishbone_bd_ram_mem3_92_25, p_wishbone_bd_ram_mem3_92_26,
         p_wishbone_bd_ram_mem3_92_27, p_wishbone_bd_ram_mem3_92_28,
         p_wishbone_bd_ram_mem3_92_29, p_wishbone_bd_ram_mem3_92_30,
         p_wishbone_bd_ram_mem3_92_31, p_wishbone_bd_ram_mem3_93_24,
         p_wishbone_bd_ram_mem3_93_25, p_wishbone_bd_ram_mem3_93_26,
         p_wishbone_bd_ram_mem3_93_27, p_wishbone_bd_ram_mem3_93_28,
         p_wishbone_bd_ram_mem3_93_29, p_wishbone_bd_ram_mem3_93_30,
         p_wishbone_bd_ram_mem3_93_31, p_wishbone_bd_ram_mem3_94_24,
         p_wishbone_bd_ram_mem3_94_25, p_wishbone_bd_ram_mem3_94_26,
         p_wishbone_bd_ram_mem3_94_27, p_wishbone_bd_ram_mem3_94_28,
         p_wishbone_bd_ram_mem3_94_29, p_wishbone_bd_ram_mem3_94_30,
         p_wishbone_bd_ram_mem3_94_31, p_wishbone_bd_ram_mem3_95_24,
         p_wishbone_bd_ram_mem3_95_25, p_wishbone_bd_ram_mem3_95_26,
         p_wishbone_bd_ram_mem3_95_27, p_wishbone_bd_ram_mem3_95_28,
         p_wishbone_bd_ram_mem3_95_29, p_wishbone_bd_ram_mem3_95_30,
         p_wishbone_bd_ram_mem3_95_31, p_wishbone_bd_ram_mem3_96_24,
         p_wishbone_bd_ram_mem3_96_25, p_wishbone_bd_ram_mem3_96_26,
         p_wishbone_bd_ram_mem3_96_27, p_wishbone_bd_ram_mem3_96_28,
         p_wishbone_bd_ram_mem3_96_29, p_wishbone_bd_ram_mem3_96_30,
         p_wishbone_bd_ram_mem3_96_31, p_wishbone_bd_ram_mem3_97_24,
         p_wishbone_bd_ram_mem3_97_25, p_wishbone_bd_ram_mem3_97_26,
         p_wishbone_bd_ram_mem3_97_27, p_wishbone_bd_ram_mem3_97_28,
         p_wishbone_bd_ram_mem3_97_29, p_wishbone_bd_ram_mem3_97_30,
         p_wishbone_bd_ram_mem3_97_31, p_wishbone_bd_ram_mem3_98_24,
         p_wishbone_bd_ram_mem3_98_25, p_wishbone_bd_ram_mem3_98_26,
         p_wishbone_bd_ram_mem3_98_27, p_wishbone_bd_ram_mem3_98_28,
         p_wishbone_bd_ram_mem3_98_29, p_wishbone_bd_ram_mem3_98_30,
         p_wishbone_bd_ram_mem3_98_31, p_wishbone_bd_ram_mem3_99_24,
         p_wishbone_bd_ram_mem3_99_25, p_wishbone_bd_ram_mem3_99_26,
         p_wishbone_bd_ram_mem3_99_27, p_wishbone_bd_ram_mem3_99_28,
         p_wishbone_bd_ram_mem3_99_29, p_wishbone_bd_ram_mem3_99_30,
         p_wishbone_bd_ram_mem3_99_31, p_wishbone_bd_ram_mem3_100_24,
         p_wishbone_bd_ram_mem3_100_25, p_wishbone_bd_ram_mem3_100_26,
         p_wishbone_bd_ram_mem3_100_27, p_wishbone_bd_ram_mem3_100_28,
         p_wishbone_bd_ram_mem3_100_29, p_wishbone_bd_ram_mem3_100_30,
         p_wishbone_bd_ram_mem3_100_31, p_wishbone_bd_ram_mem3_101_24,
         p_wishbone_bd_ram_mem3_101_25, p_wishbone_bd_ram_mem3_101_26,
         p_wishbone_bd_ram_mem3_101_27, p_wishbone_bd_ram_mem3_101_28,
         p_wishbone_bd_ram_mem3_101_29, p_wishbone_bd_ram_mem3_101_30,
         p_wishbone_bd_ram_mem3_101_31, p_wishbone_bd_ram_mem3_102_24,
         p_wishbone_bd_ram_mem3_102_25, p_wishbone_bd_ram_mem3_102_26,
         p_wishbone_bd_ram_mem3_102_27, p_wishbone_bd_ram_mem3_102_28,
         p_wishbone_bd_ram_mem3_102_29, p_wishbone_bd_ram_mem3_102_30,
         p_wishbone_bd_ram_mem3_102_31, p_wishbone_bd_ram_mem3_103_24,
         p_wishbone_bd_ram_mem3_103_25, p_wishbone_bd_ram_mem3_103_26,
         p_wishbone_bd_ram_mem3_103_27, p_wishbone_bd_ram_mem3_103_28,
         p_wishbone_bd_ram_mem3_103_29, p_wishbone_bd_ram_mem3_103_30,
         p_wishbone_bd_ram_mem3_103_31, p_wishbone_bd_ram_mem3_104_24,
         p_wishbone_bd_ram_mem3_104_25, p_wishbone_bd_ram_mem3_104_26,
         p_wishbone_bd_ram_mem3_104_27, p_wishbone_bd_ram_mem3_104_28,
         p_wishbone_bd_ram_mem3_104_29, p_wishbone_bd_ram_mem3_104_30,
         p_wishbone_bd_ram_mem3_104_31, p_wishbone_bd_ram_mem3_105_24,
         p_wishbone_bd_ram_mem3_105_25, p_wishbone_bd_ram_mem3_105_26,
         p_wishbone_bd_ram_mem3_105_27, p_wishbone_bd_ram_mem3_105_28,
         p_wishbone_bd_ram_mem3_105_29, p_wishbone_bd_ram_mem3_105_30,
         p_wishbone_bd_ram_mem3_105_31, p_wishbone_bd_ram_mem3_106_24,
         p_wishbone_bd_ram_mem3_106_25, p_wishbone_bd_ram_mem3_106_26,
         p_wishbone_bd_ram_mem3_106_27, p_wishbone_bd_ram_mem3_106_28,
         p_wishbone_bd_ram_mem3_106_29, p_wishbone_bd_ram_mem3_106_30,
         p_wishbone_bd_ram_mem3_106_31, p_wishbone_bd_ram_mem3_107_24,
         p_wishbone_bd_ram_mem3_107_25, p_wishbone_bd_ram_mem3_107_26,
         p_wishbone_bd_ram_mem3_107_27, p_wishbone_bd_ram_mem3_107_28,
         p_wishbone_bd_ram_mem3_107_29, p_wishbone_bd_ram_mem3_107_30,
         p_wishbone_bd_ram_mem3_107_31, p_wishbone_bd_ram_mem3_108_24,
         p_wishbone_bd_ram_mem3_108_25, p_wishbone_bd_ram_mem3_108_26,
         p_wishbone_bd_ram_mem3_108_27, p_wishbone_bd_ram_mem3_108_28,
         p_wishbone_bd_ram_mem3_108_29, p_wishbone_bd_ram_mem3_108_30,
         p_wishbone_bd_ram_mem3_108_31, p_wishbone_bd_ram_mem3_109_24,
         p_wishbone_bd_ram_mem3_109_25, p_wishbone_bd_ram_mem3_109_26,
         p_wishbone_bd_ram_mem3_109_27, p_wishbone_bd_ram_mem3_109_28,
         p_wishbone_bd_ram_mem3_109_29, p_wishbone_bd_ram_mem3_109_30,
         p_wishbone_bd_ram_mem3_109_31, p_wishbone_bd_ram_mem3_110_24,
         p_wishbone_bd_ram_mem3_110_25, p_wishbone_bd_ram_mem3_110_26,
         p_wishbone_bd_ram_mem3_110_27, p_wishbone_bd_ram_mem3_110_28,
         p_wishbone_bd_ram_mem3_110_29, p_wishbone_bd_ram_mem3_110_30,
         p_wishbone_bd_ram_mem3_110_31, p_wishbone_bd_ram_mem3_111_24,
         p_wishbone_bd_ram_mem3_111_25, p_wishbone_bd_ram_mem3_111_26,
         p_wishbone_bd_ram_mem3_111_27, p_wishbone_bd_ram_mem3_111_28,
         p_wishbone_bd_ram_mem3_111_29, p_wishbone_bd_ram_mem3_111_30,
         p_wishbone_bd_ram_mem3_111_31, p_wishbone_bd_ram_mem3_112_24,
         p_wishbone_bd_ram_mem3_112_25, p_wishbone_bd_ram_mem3_112_26,
         p_wishbone_bd_ram_mem3_112_27, p_wishbone_bd_ram_mem3_112_28,
         p_wishbone_bd_ram_mem3_112_29, p_wishbone_bd_ram_mem3_112_30,
         p_wishbone_bd_ram_mem3_112_31, p_wishbone_bd_ram_mem3_113_24,
         p_wishbone_bd_ram_mem3_113_25, p_wishbone_bd_ram_mem3_113_26,
         p_wishbone_bd_ram_mem3_113_27, p_wishbone_bd_ram_mem3_113_28,
         p_wishbone_bd_ram_mem3_113_29, p_wishbone_bd_ram_mem3_113_30,
         p_wishbone_bd_ram_mem3_113_31, p_wishbone_bd_ram_mem3_114_24,
         p_wishbone_bd_ram_mem3_114_25, p_wishbone_bd_ram_mem3_114_26,
         p_wishbone_bd_ram_mem3_114_27, p_wishbone_bd_ram_mem3_114_28,
         p_wishbone_bd_ram_mem3_114_29, p_wishbone_bd_ram_mem3_114_30,
         p_wishbone_bd_ram_mem3_114_31, p_wishbone_bd_ram_mem3_115_24,
         p_wishbone_bd_ram_mem3_115_25, p_wishbone_bd_ram_mem3_115_26,
         p_wishbone_bd_ram_mem3_115_27, p_wishbone_bd_ram_mem3_115_28,
         p_wishbone_bd_ram_mem3_115_29, p_wishbone_bd_ram_mem3_115_30,
         p_wishbone_bd_ram_mem3_115_31, p_wishbone_bd_ram_mem3_116_24,
         p_wishbone_bd_ram_mem3_116_25, p_wishbone_bd_ram_mem3_116_26,
         p_wishbone_bd_ram_mem3_116_27, p_wishbone_bd_ram_mem3_116_28,
         p_wishbone_bd_ram_mem3_116_29, p_wishbone_bd_ram_mem3_116_30,
         p_wishbone_bd_ram_mem3_116_31, p_wishbone_bd_ram_mem3_117_24,
         p_wishbone_bd_ram_mem3_117_25, p_wishbone_bd_ram_mem3_117_26,
         p_wishbone_bd_ram_mem3_117_27, p_wishbone_bd_ram_mem3_117_28,
         p_wishbone_bd_ram_mem3_117_29, p_wishbone_bd_ram_mem3_117_30,
         p_wishbone_bd_ram_mem3_117_31, p_wishbone_bd_ram_mem3_118_24,
         p_wishbone_bd_ram_mem3_118_25, p_wishbone_bd_ram_mem3_118_26,
         p_wishbone_bd_ram_mem3_118_27, p_wishbone_bd_ram_mem3_118_28,
         p_wishbone_bd_ram_mem3_118_29, p_wishbone_bd_ram_mem3_118_30,
         p_wishbone_bd_ram_mem3_118_31, p_wishbone_bd_ram_mem3_119_24,
         p_wishbone_bd_ram_mem3_119_25, p_wishbone_bd_ram_mem3_119_26,
         p_wishbone_bd_ram_mem3_119_27, p_wishbone_bd_ram_mem3_119_28,
         p_wishbone_bd_ram_mem3_119_29, p_wishbone_bd_ram_mem3_119_30,
         p_wishbone_bd_ram_mem3_119_31, p_wishbone_bd_ram_mem3_120_24,
         p_wishbone_bd_ram_mem3_120_25, p_wishbone_bd_ram_mem3_120_26,
         p_wishbone_bd_ram_mem3_120_27, p_wishbone_bd_ram_mem3_120_28,
         p_wishbone_bd_ram_mem3_120_29, p_wishbone_bd_ram_mem3_120_30,
         p_wishbone_bd_ram_mem3_120_31, p_wishbone_bd_ram_mem3_121_24,
         p_wishbone_bd_ram_mem3_121_25, p_wishbone_bd_ram_mem3_121_26,
         p_wishbone_bd_ram_mem3_121_27, p_wishbone_bd_ram_mem3_121_28,
         p_wishbone_bd_ram_mem3_121_29, p_wishbone_bd_ram_mem3_121_30,
         p_wishbone_bd_ram_mem3_121_31, p_wishbone_bd_ram_mem3_122_24,
         p_wishbone_bd_ram_mem3_122_25, p_wishbone_bd_ram_mem3_122_26,
         p_wishbone_bd_ram_mem3_122_27, p_wishbone_bd_ram_mem3_122_28,
         p_wishbone_bd_ram_mem3_122_29, p_wishbone_bd_ram_mem3_122_30,
         p_wishbone_bd_ram_mem3_122_31, p_wishbone_bd_ram_mem3_123_24,
         p_wishbone_bd_ram_mem3_123_25, p_wishbone_bd_ram_mem3_123_26,
         p_wishbone_bd_ram_mem3_123_27, p_wishbone_bd_ram_mem3_123_28,
         p_wishbone_bd_ram_mem3_123_29, p_wishbone_bd_ram_mem3_123_30,
         p_wishbone_bd_ram_mem3_123_31, p_wishbone_bd_ram_mem3_124_24,
         p_wishbone_bd_ram_mem3_124_25, p_wishbone_bd_ram_mem3_124_26,
         p_wishbone_bd_ram_mem3_124_27, p_wishbone_bd_ram_mem3_124_28,
         p_wishbone_bd_ram_mem3_124_29, p_wishbone_bd_ram_mem3_124_30,
         p_wishbone_bd_ram_mem3_124_31, p_wishbone_bd_ram_mem3_125_24,
         p_wishbone_bd_ram_mem3_125_25, p_wishbone_bd_ram_mem3_125_26,
         p_wishbone_bd_ram_mem3_125_27, p_wishbone_bd_ram_mem3_125_28,
         p_wishbone_bd_ram_mem3_125_29, p_wishbone_bd_ram_mem3_125_30,
         p_wishbone_bd_ram_mem3_125_31, p_wishbone_bd_ram_mem3_126_24,
         p_wishbone_bd_ram_mem3_126_25, p_wishbone_bd_ram_mem3_126_26,
         p_wishbone_bd_ram_mem3_126_27, p_wishbone_bd_ram_mem3_126_28,
         p_wishbone_bd_ram_mem3_126_29, p_wishbone_bd_ram_mem3_126_30,
         p_wishbone_bd_ram_mem3_126_31, p_wishbone_bd_ram_mem3_127_24,
         p_wishbone_bd_ram_mem3_127_25, p_wishbone_bd_ram_mem3_127_26,
         p_wishbone_bd_ram_mem3_127_27, p_wishbone_bd_ram_mem3_127_28,
         p_wishbone_bd_ram_mem3_127_29, p_wishbone_bd_ram_mem3_127_30,
         p_wishbone_bd_ram_mem3_127_31, p_wishbone_bd_ram_mem3_128_24,
         p_wishbone_bd_ram_mem3_128_25, p_wishbone_bd_ram_mem3_128_26,
         p_wishbone_bd_ram_mem3_128_27, p_wishbone_bd_ram_mem3_128_28,
         p_wishbone_bd_ram_mem3_128_29, p_wishbone_bd_ram_mem3_128_30,
         p_wishbone_bd_ram_mem3_128_31, p_wishbone_bd_ram_mem3_129_24,
         p_wishbone_bd_ram_mem3_129_25, p_wishbone_bd_ram_mem3_129_26,
         p_wishbone_bd_ram_mem3_129_27, p_wishbone_bd_ram_mem3_129_28,
         p_wishbone_bd_ram_mem3_129_29, p_wishbone_bd_ram_mem3_129_30,
         p_wishbone_bd_ram_mem3_129_31, p_wishbone_bd_ram_mem3_130_24,
         p_wishbone_bd_ram_mem3_130_25, p_wishbone_bd_ram_mem3_130_26,
         p_wishbone_bd_ram_mem3_130_27, p_wishbone_bd_ram_mem3_130_28,
         p_wishbone_bd_ram_mem3_130_29, p_wishbone_bd_ram_mem3_130_30,
         p_wishbone_bd_ram_mem3_130_31, p_wishbone_bd_ram_mem3_131_24,
         p_wishbone_bd_ram_mem3_131_25, p_wishbone_bd_ram_mem3_131_26,
         p_wishbone_bd_ram_mem3_131_27, p_wishbone_bd_ram_mem3_131_28,
         p_wishbone_bd_ram_mem3_131_29, p_wishbone_bd_ram_mem3_131_30,
         p_wishbone_bd_ram_mem3_131_31, p_wishbone_bd_ram_mem3_132_24,
         p_wishbone_bd_ram_mem3_132_25, p_wishbone_bd_ram_mem3_132_26,
         p_wishbone_bd_ram_mem3_132_27, p_wishbone_bd_ram_mem3_132_28,
         p_wishbone_bd_ram_mem3_132_29, p_wishbone_bd_ram_mem3_132_30,
         p_wishbone_bd_ram_mem3_132_31, p_wishbone_bd_ram_mem3_133_24,
         p_wishbone_bd_ram_mem3_133_25, p_wishbone_bd_ram_mem3_133_26,
         p_wishbone_bd_ram_mem3_133_27, p_wishbone_bd_ram_mem3_133_28,
         p_wishbone_bd_ram_mem3_133_29, p_wishbone_bd_ram_mem3_133_30,
         p_wishbone_bd_ram_mem3_133_31, p_wishbone_bd_ram_mem3_134_24,
         p_wishbone_bd_ram_mem3_134_25, p_wishbone_bd_ram_mem3_134_26,
         p_wishbone_bd_ram_mem3_134_27, p_wishbone_bd_ram_mem3_134_28,
         p_wishbone_bd_ram_mem3_134_29, p_wishbone_bd_ram_mem3_134_30,
         p_wishbone_bd_ram_mem3_134_31, p_wishbone_bd_ram_mem3_135_24,
         p_wishbone_bd_ram_mem3_135_25, p_wishbone_bd_ram_mem3_135_26,
         p_wishbone_bd_ram_mem3_135_27, p_wishbone_bd_ram_mem3_135_28,
         p_wishbone_bd_ram_mem3_135_29, p_wishbone_bd_ram_mem3_135_30,
         p_wishbone_bd_ram_mem3_135_31, p_wishbone_bd_ram_mem3_136_24,
         p_wishbone_bd_ram_mem3_136_25, p_wishbone_bd_ram_mem3_136_26,
         p_wishbone_bd_ram_mem3_136_27, p_wishbone_bd_ram_mem3_136_28,
         p_wishbone_bd_ram_mem3_136_29, p_wishbone_bd_ram_mem3_136_30,
         p_wishbone_bd_ram_mem3_136_31, p_wishbone_bd_ram_mem3_137_24,
         p_wishbone_bd_ram_mem3_137_25, p_wishbone_bd_ram_mem3_137_26,
         p_wishbone_bd_ram_mem3_137_27, p_wishbone_bd_ram_mem3_137_28,
         p_wishbone_bd_ram_mem3_137_29, p_wishbone_bd_ram_mem3_137_30,
         p_wishbone_bd_ram_mem3_137_31, p_wishbone_bd_ram_mem3_138_24,
         p_wishbone_bd_ram_mem3_138_25, p_wishbone_bd_ram_mem3_138_26,
         p_wishbone_bd_ram_mem3_138_27, p_wishbone_bd_ram_mem3_138_28,
         p_wishbone_bd_ram_mem3_138_29, p_wishbone_bd_ram_mem3_138_30,
         p_wishbone_bd_ram_mem3_138_31, p_wishbone_bd_ram_mem3_139_24,
         p_wishbone_bd_ram_mem3_139_25, p_wishbone_bd_ram_mem3_139_26,
         p_wishbone_bd_ram_mem3_139_27, p_wishbone_bd_ram_mem3_139_28,
         p_wishbone_bd_ram_mem3_139_29, p_wishbone_bd_ram_mem3_139_30,
         p_wishbone_bd_ram_mem3_139_31, p_wishbone_bd_ram_mem3_140_24,
         p_wishbone_bd_ram_mem3_140_25, p_wishbone_bd_ram_mem3_140_26,
         p_wishbone_bd_ram_mem3_140_27, p_wishbone_bd_ram_mem3_140_28,
         p_wishbone_bd_ram_mem3_140_29, p_wishbone_bd_ram_mem3_140_30,
         p_wishbone_bd_ram_mem3_140_31, p_wishbone_bd_ram_mem3_141_24,
         p_wishbone_bd_ram_mem3_141_25, p_wishbone_bd_ram_mem3_141_26,
         p_wishbone_bd_ram_mem3_141_27, p_wishbone_bd_ram_mem3_141_28,
         p_wishbone_bd_ram_mem3_141_29, p_wishbone_bd_ram_mem3_141_30,
         p_wishbone_bd_ram_mem3_141_31, p_wishbone_bd_ram_mem3_142_24,
         p_wishbone_bd_ram_mem3_142_25, p_wishbone_bd_ram_mem3_142_26,
         p_wishbone_bd_ram_mem3_142_27, p_wishbone_bd_ram_mem3_142_28,
         p_wishbone_bd_ram_mem3_142_29, p_wishbone_bd_ram_mem3_142_30,
         p_wishbone_bd_ram_mem3_142_31, p_wishbone_bd_ram_mem3_143_24,
         p_wishbone_bd_ram_mem3_143_25, p_wishbone_bd_ram_mem3_143_26,
         p_wishbone_bd_ram_mem3_143_27, p_wishbone_bd_ram_mem3_143_28,
         p_wishbone_bd_ram_mem3_143_29, p_wishbone_bd_ram_mem3_143_30,
         p_wishbone_bd_ram_mem3_143_31, p_wishbone_bd_ram_mem3_144_24,
         p_wishbone_bd_ram_mem3_144_25, p_wishbone_bd_ram_mem3_144_26,
         p_wishbone_bd_ram_mem3_144_27, p_wishbone_bd_ram_mem3_144_28,
         p_wishbone_bd_ram_mem3_144_29, p_wishbone_bd_ram_mem3_144_30,
         p_wishbone_bd_ram_mem3_144_31, p_wishbone_bd_ram_mem3_145_24,
         p_wishbone_bd_ram_mem3_145_25, p_wishbone_bd_ram_mem3_145_26,
         p_wishbone_bd_ram_mem3_145_27, p_wishbone_bd_ram_mem3_145_28,
         p_wishbone_bd_ram_mem3_145_29, p_wishbone_bd_ram_mem3_145_30,
         p_wishbone_bd_ram_mem3_145_31, p_wishbone_bd_ram_mem3_146_24,
         p_wishbone_bd_ram_mem3_146_25, p_wishbone_bd_ram_mem3_146_26,
         p_wishbone_bd_ram_mem3_146_27, p_wishbone_bd_ram_mem3_146_28,
         p_wishbone_bd_ram_mem3_146_29, p_wishbone_bd_ram_mem3_146_30,
         p_wishbone_bd_ram_mem3_146_31, p_wishbone_bd_ram_mem3_147_24,
         p_wishbone_bd_ram_mem3_147_25, p_wishbone_bd_ram_mem3_147_26,
         p_wishbone_bd_ram_mem3_147_27, p_wishbone_bd_ram_mem3_147_28,
         p_wishbone_bd_ram_mem3_147_29, p_wishbone_bd_ram_mem3_147_30,
         p_wishbone_bd_ram_mem3_147_31, p_wishbone_bd_ram_mem3_148_24,
         p_wishbone_bd_ram_mem3_148_25, p_wishbone_bd_ram_mem3_148_26,
         p_wishbone_bd_ram_mem3_148_27, p_wishbone_bd_ram_mem3_148_28,
         p_wishbone_bd_ram_mem3_148_29, p_wishbone_bd_ram_mem3_148_30,
         p_wishbone_bd_ram_mem3_148_31, p_wishbone_bd_ram_mem3_149_24,
         p_wishbone_bd_ram_mem3_149_25, p_wishbone_bd_ram_mem3_149_26,
         p_wishbone_bd_ram_mem3_149_27, p_wishbone_bd_ram_mem3_149_28,
         p_wishbone_bd_ram_mem3_149_29, p_wishbone_bd_ram_mem3_149_30,
         p_wishbone_bd_ram_mem3_149_31, p_wishbone_bd_ram_mem3_150_24,
         p_wishbone_bd_ram_mem3_150_25, p_wishbone_bd_ram_mem3_150_26,
         p_wishbone_bd_ram_mem3_150_27, p_wishbone_bd_ram_mem3_150_28,
         p_wishbone_bd_ram_mem3_150_29, p_wishbone_bd_ram_mem3_150_30,
         p_wishbone_bd_ram_mem3_150_31, p_wishbone_bd_ram_mem3_151_24,
         p_wishbone_bd_ram_mem3_151_25, p_wishbone_bd_ram_mem3_151_26,
         p_wishbone_bd_ram_mem3_151_27, p_wishbone_bd_ram_mem3_151_28,
         p_wishbone_bd_ram_mem3_151_29, p_wishbone_bd_ram_mem3_151_30,
         p_wishbone_bd_ram_mem3_151_31, p_wishbone_bd_ram_mem3_152_24,
         p_wishbone_bd_ram_mem3_152_25, p_wishbone_bd_ram_mem3_152_26,
         p_wishbone_bd_ram_mem3_152_27, p_wishbone_bd_ram_mem3_152_28,
         p_wishbone_bd_ram_mem3_152_29, p_wishbone_bd_ram_mem3_152_30,
         p_wishbone_bd_ram_mem3_152_31, p_wishbone_bd_ram_mem3_153_24,
         p_wishbone_bd_ram_mem3_153_25, p_wishbone_bd_ram_mem3_153_26,
         p_wishbone_bd_ram_mem3_153_27, p_wishbone_bd_ram_mem3_153_28,
         p_wishbone_bd_ram_mem3_153_29, p_wishbone_bd_ram_mem3_153_30,
         p_wishbone_bd_ram_mem3_153_31, p_wishbone_bd_ram_mem3_154_24,
         p_wishbone_bd_ram_mem3_154_25, p_wishbone_bd_ram_mem3_154_26,
         p_wishbone_bd_ram_mem3_154_27, p_wishbone_bd_ram_mem3_154_28,
         p_wishbone_bd_ram_mem3_154_29, p_wishbone_bd_ram_mem3_154_30,
         p_wishbone_bd_ram_mem3_154_31, p_wishbone_bd_ram_mem3_155_24,
         p_wishbone_bd_ram_mem3_155_25, p_wishbone_bd_ram_mem3_155_26,
         p_wishbone_bd_ram_mem3_155_27, p_wishbone_bd_ram_mem3_155_28,
         p_wishbone_bd_ram_mem3_155_29, p_wishbone_bd_ram_mem3_155_30,
         p_wishbone_bd_ram_mem3_155_31, p_wishbone_bd_ram_mem3_156_24,
         p_wishbone_bd_ram_mem3_156_25, p_wishbone_bd_ram_mem3_156_26,
         p_wishbone_bd_ram_mem3_156_27, p_wishbone_bd_ram_mem3_156_28,
         p_wishbone_bd_ram_mem3_156_29, p_wishbone_bd_ram_mem3_156_30,
         p_wishbone_bd_ram_mem3_156_31, p_wishbone_bd_ram_mem3_157_24,
         p_wishbone_bd_ram_mem3_157_25, p_wishbone_bd_ram_mem3_157_26,
         p_wishbone_bd_ram_mem3_157_27, p_wishbone_bd_ram_mem3_157_28,
         p_wishbone_bd_ram_mem3_157_29, p_wishbone_bd_ram_mem3_157_30,
         p_wishbone_bd_ram_mem3_157_31, p_wishbone_bd_ram_mem3_158_24,
         p_wishbone_bd_ram_mem3_158_25, p_wishbone_bd_ram_mem3_158_26,
         p_wishbone_bd_ram_mem3_158_27, p_wishbone_bd_ram_mem3_158_28,
         p_wishbone_bd_ram_mem3_158_29, p_wishbone_bd_ram_mem3_158_30,
         p_wishbone_bd_ram_mem3_158_31, p_wishbone_bd_ram_mem3_159_24,
         p_wishbone_bd_ram_mem3_159_25, p_wishbone_bd_ram_mem3_159_26,
         p_wishbone_bd_ram_mem3_159_27, p_wishbone_bd_ram_mem3_159_28,
         p_wishbone_bd_ram_mem3_159_29, p_wishbone_bd_ram_mem3_159_30,
         p_wishbone_bd_ram_mem3_159_31, p_wishbone_bd_ram_mem3_160_24,
         p_wishbone_bd_ram_mem3_160_25, p_wishbone_bd_ram_mem3_160_26,
         p_wishbone_bd_ram_mem3_160_27, p_wishbone_bd_ram_mem3_160_28,
         p_wishbone_bd_ram_mem3_160_29, p_wishbone_bd_ram_mem3_160_30,
         p_wishbone_bd_ram_mem3_160_31, p_wishbone_bd_ram_mem3_161_24,
         p_wishbone_bd_ram_mem3_161_25, p_wishbone_bd_ram_mem3_161_26,
         p_wishbone_bd_ram_mem3_161_27, p_wishbone_bd_ram_mem3_161_28,
         p_wishbone_bd_ram_mem3_161_29, p_wishbone_bd_ram_mem3_161_30,
         p_wishbone_bd_ram_mem3_161_31, p_wishbone_bd_ram_mem3_162_24,
         p_wishbone_bd_ram_mem3_162_25, p_wishbone_bd_ram_mem3_162_26,
         p_wishbone_bd_ram_mem3_162_27, p_wishbone_bd_ram_mem3_162_28,
         p_wishbone_bd_ram_mem3_162_29, p_wishbone_bd_ram_mem3_162_30,
         p_wishbone_bd_ram_mem3_162_31, p_wishbone_bd_ram_mem3_163_24,
         p_wishbone_bd_ram_mem3_163_25, p_wishbone_bd_ram_mem3_163_26,
         p_wishbone_bd_ram_mem3_163_27, p_wishbone_bd_ram_mem3_163_28,
         p_wishbone_bd_ram_mem3_163_29, p_wishbone_bd_ram_mem3_163_30,
         p_wishbone_bd_ram_mem3_163_31, p_wishbone_bd_ram_mem3_164_24,
         p_wishbone_bd_ram_mem3_164_25, p_wishbone_bd_ram_mem3_164_26,
         p_wishbone_bd_ram_mem3_164_27, p_wishbone_bd_ram_mem3_164_28,
         p_wishbone_bd_ram_mem3_164_29, p_wishbone_bd_ram_mem3_164_30,
         p_wishbone_bd_ram_mem3_164_31, p_wishbone_bd_ram_mem3_165_24,
         p_wishbone_bd_ram_mem3_165_25, p_wishbone_bd_ram_mem3_165_26,
         p_wishbone_bd_ram_mem3_165_27, p_wishbone_bd_ram_mem3_165_28,
         p_wishbone_bd_ram_mem3_165_29, p_wishbone_bd_ram_mem3_165_30,
         p_wishbone_bd_ram_mem3_165_31, p_wishbone_bd_ram_mem3_166_24,
         p_wishbone_bd_ram_mem3_166_25, p_wishbone_bd_ram_mem3_166_26,
         p_wishbone_bd_ram_mem3_166_27, p_wishbone_bd_ram_mem3_166_28,
         p_wishbone_bd_ram_mem3_166_29, p_wishbone_bd_ram_mem3_166_30,
         p_wishbone_bd_ram_mem3_166_31, p_wishbone_bd_ram_mem3_167_24,
         p_wishbone_bd_ram_mem3_167_25, p_wishbone_bd_ram_mem3_167_26,
         p_wishbone_bd_ram_mem3_167_27, p_wishbone_bd_ram_mem3_167_28,
         p_wishbone_bd_ram_mem3_167_29, p_wishbone_bd_ram_mem3_167_30,
         p_wishbone_bd_ram_mem3_167_31, p_wishbone_bd_ram_mem3_168_24,
         p_wishbone_bd_ram_mem3_168_25, p_wishbone_bd_ram_mem3_168_26,
         p_wishbone_bd_ram_mem3_168_27, p_wishbone_bd_ram_mem3_168_28,
         p_wishbone_bd_ram_mem3_168_29, p_wishbone_bd_ram_mem3_168_30,
         p_wishbone_bd_ram_mem3_168_31, p_wishbone_bd_ram_mem3_169_24,
         p_wishbone_bd_ram_mem3_169_25, p_wishbone_bd_ram_mem3_169_26,
         p_wishbone_bd_ram_mem3_169_27, p_wishbone_bd_ram_mem3_169_28,
         p_wishbone_bd_ram_mem3_169_29, p_wishbone_bd_ram_mem3_169_30,
         p_wishbone_bd_ram_mem3_169_31, p_wishbone_bd_ram_mem3_170_24,
         p_wishbone_bd_ram_mem3_170_25, p_wishbone_bd_ram_mem3_170_26,
         p_wishbone_bd_ram_mem3_170_27, p_wishbone_bd_ram_mem3_170_28,
         p_wishbone_bd_ram_mem3_170_29, p_wishbone_bd_ram_mem3_170_30,
         p_wishbone_bd_ram_mem3_170_31, p_wishbone_bd_ram_mem3_171_24,
         p_wishbone_bd_ram_mem3_171_25, p_wishbone_bd_ram_mem3_171_26,
         p_wishbone_bd_ram_mem3_171_27, p_wishbone_bd_ram_mem3_171_28,
         p_wishbone_bd_ram_mem3_171_29, p_wishbone_bd_ram_mem3_171_30,
         p_wishbone_bd_ram_mem3_171_31, p_wishbone_bd_ram_mem3_172_24,
         p_wishbone_bd_ram_mem3_172_25, p_wishbone_bd_ram_mem3_172_26,
         p_wishbone_bd_ram_mem3_172_27, p_wishbone_bd_ram_mem3_172_28,
         p_wishbone_bd_ram_mem3_172_29, p_wishbone_bd_ram_mem3_172_30,
         p_wishbone_bd_ram_mem3_172_31, p_wishbone_bd_ram_mem3_173_24,
         p_wishbone_bd_ram_mem3_173_25, p_wishbone_bd_ram_mem3_173_26,
         p_wishbone_bd_ram_mem3_173_27, p_wishbone_bd_ram_mem3_173_28,
         p_wishbone_bd_ram_mem3_173_29, p_wishbone_bd_ram_mem3_173_30,
         p_wishbone_bd_ram_mem3_173_31, p_wishbone_bd_ram_mem3_174_24,
         p_wishbone_bd_ram_mem3_174_25, p_wishbone_bd_ram_mem3_174_26,
         p_wishbone_bd_ram_mem3_174_27, p_wishbone_bd_ram_mem3_174_28,
         p_wishbone_bd_ram_mem3_174_29, p_wishbone_bd_ram_mem3_174_30,
         p_wishbone_bd_ram_mem3_174_31, p_wishbone_bd_ram_mem3_175_24,
         p_wishbone_bd_ram_mem3_175_25, p_wishbone_bd_ram_mem3_175_26,
         p_wishbone_bd_ram_mem3_175_27, p_wishbone_bd_ram_mem3_175_28,
         p_wishbone_bd_ram_mem3_175_29, p_wishbone_bd_ram_mem3_175_30,
         p_wishbone_bd_ram_mem3_175_31, p_wishbone_bd_ram_mem3_176_24,
         p_wishbone_bd_ram_mem3_176_25, p_wishbone_bd_ram_mem3_176_26,
         p_wishbone_bd_ram_mem3_176_27, p_wishbone_bd_ram_mem3_176_28,
         p_wishbone_bd_ram_mem3_176_29, p_wishbone_bd_ram_mem3_176_30,
         p_wishbone_bd_ram_mem3_176_31, p_wishbone_bd_ram_mem3_177_24,
         p_wishbone_bd_ram_mem3_177_25, p_wishbone_bd_ram_mem3_177_26,
         p_wishbone_bd_ram_mem3_177_27, p_wishbone_bd_ram_mem3_177_28,
         p_wishbone_bd_ram_mem3_177_29, p_wishbone_bd_ram_mem3_177_30,
         p_wishbone_bd_ram_mem3_177_31, p_wishbone_bd_ram_mem3_178_24,
         p_wishbone_bd_ram_mem3_178_25, p_wishbone_bd_ram_mem3_178_26,
         p_wishbone_bd_ram_mem3_178_27, p_wishbone_bd_ram_mem3_178_28,
         p_wishbone_bd_ram_mem3_178_29, p_wishbone_bd_ram_mem3_178_30,
         p_wishbone_bd_ram_mem3_178_31, p_wishbone_bd_ram_mem3_179_24,
         p_wishbone_bd_ram_mem3_179_25, p_wishbone_bd_ram_mem3_179_26,
         p_wishbone_bd_ram_mem3_179_27, p_wishbone_bd_ram_mem3_179_28,
         p_wishbone_bd_ram_mem3_179_29, p_wishbone_bd_ram_mem3_179_30,
         p_wishbone_bd_ram_mem3_179_31, p_wishbone_bd_ram_mem3_180_24,
         p_wishbone_bd_ram_mem3_180_25, p_wishbone_bd_ram_mem3_180_26,
         p_wishbone_bd_ram_mem3_180_27, p_wishbone_bd_ram_mem3_180_28,
         p_wishbone_bd_ram_mem3_180_29, p_wishbone_bd_ram_mem3_180_30,
         p_wishbone_bd_ram_mem3_180_31, p_wishbone_bd_ram_mem3_181_24,
         p_wishbone_bd_ram_mem3_181_25, p_wishbone_bd_ram_mem3_181_26,
         p_wishbone_bd_ram_mem3_181_27, p_wishbone_bd_ram_mem3_181_28,
         p_wishbone_bd_ram_mem3_181_29, p_wishbone_bd_ram_mem3_181_30,
         p_wishbone_bd_ram_mem3_181_31, p_wishbone_bd_ram_mem3_182_24,
         p_wishbone_bd_ram_mem3_182_25, p_wishbone_bd_ram_mem3_182_26,
         p_wishbone_bd_ram_mem3_182_27, p_wishbone_bd_ram_mem3_182_28,
         p_wishbone_bd_ram_mem3_182_29, p_wishbone_bd_ram_mem3_182_30,
         p_wishbone_bd_ram_mem3_182_31, p_wishbone_bd_ram_mem3_183_24,
         p_wishbone_bd_ram_mem3_183_25, p_wishbone_bd_ram_mem3_183_26,
         p_wishbone_bd_ram_mem3_183_27, p_wishbone_bd_ram_mem3_183_28,
         p_wishbone_bd_ram_mem3_183_29, p_wishbone_bd_ram_mem3_183_30,
         p_wishbone_bd_ram_mem3_183_31, p_wishbone_bd_ram_mem3_184_24,
         p_wishbone_bd_ram_mem3_184_25, p_wishbone_bd_ram_mem3_184_26,
         p_wishbone_bd_ram_mem3_184_27, p_wishbone_bd_ram_mem3_184_28,
         p_wishbone_bd_ram_mem3_184_29, p_wishbone_bd_ram_mem3_184_30,
         p_wishbone_bd_ram_mem3_184_31, p_wishbone_bd_ram_mem3_185_24,
         p_wishbone_bd_ram_mem3_185_25, p_wishbone_bd_ram_mem3_185_26,
         p_wishbone_bd_ram_mem3_185_27, p_wishbone_bd_ram_mem3_185_28,
         p_wishbone_bd_ram_mem3_185_29, p_wishbone_bd_ram_mem3_185_30,
         p_wishbone_bd_ram_mem3_185_31, p_wishbone_bd_ram_mem3_186_24,
         p_wishbone_bd_ram_mem3_186_25, p_wishbone_bd_ram_mem3_186_26,
         p_wishbone_bd_ram_mem3_186_27, p_wishbone_bd_ram_mem3_186_28,
         p_wishbone_bd_ram_mem3_186_29, p_wishbone_bd_ram_mem3_186_30,
         p_wishbone_bd_ram_mem3_186_31, p_wishbone_bd_ram_mem3_187_24,
         p_wishbone_bd_ram_mem3_187_25, p_wishbone_bd_ram_mem3_187_26,
         p_wishbone_bd_ram_mem3_187_27, p_wishbone_bd_ram_mem3_187_28,
         p_wishbone_bd_ram_mem3_187_29, p_wishbone_bd_ram_mem3_187_30,
         p_wishbone_bd_ram_mem3_187_31, p_wishbone_bd_ram_mem3_188_24,
         p_wishbone_bd_ram_mem3_188_25, p_wishbone_bd_ram_mem3_188_26,
         p_wishbone_bd_ram_mem3_188_27, p_wishbone_bd_ram_mem3_188_28,
         p_wishbone_bd_ram_mem3_188_29, p_wishbone_bd_ram_mem3_188_30,
         p_wishbone_bd_ram_mem3_188_31, p_wishbone_bd_ram_mem3_189_24,
         p_wishbone_bd_ram_mem3_189_25, p_wishbone_bd_ram_mem3_189_26,
         p_wishbone_bd_ram_mem3_189_27, p_wishbone_bd_ram_mem3_189_28,
         p_wishbone_bd_ram_mem3_189_29, p_wishbone_bd_ram_mem3_189_30,
         p_wishbone_bd_ram_mem3_189_31, p_wishbone_bd_ram_mem3_190_24,
         p_wishbone_bd_ram_mem3_190_25, p_wishbone_bd_ram_mem3_190_26,
         p_wishbone_bd_ram_mem3_190_27, p_wishbone_bd_ram_mem3_190_28,
         p_wishbone_bd_ram_mem3_190_29, p_wishbone_bd_ram_mem3_190_30,
         p_wishbone_bd_ram_mem3_190_31, p_wishbone_bd_ram_mem3_191_24,
         p_wishbone_bd_ram_mem3_191_25, p_wishbone_bd_ram_mem3_191_26,
         p_wishbone_bd_ram_mem3_191_27, p_wishbone_bd_ram_mem3_191_28,
         p_wishbone_bd_ram_mem3_191_29, p_wishbone_bd_ram_mem3_191_30,
         p_wishbone_bd_ram_mem3_191_31, p_wishbone_bd_ram_mem3_192_24,
         p_wishbone_bd_ram_mem3_192_25, p_wishbone_bd_ram_mem3_192_26,
         p_wishbone_bd_ram_mem3_192_27, p_wishbone_bd_ram_mem3_192_28,
         p_wishbone_bd_ram_mem3_192_29, p_wishbone_bd_ram_mem3_192_30,
         p_wishbone_bd_ram_mem3_192_31, p_wishbone_bd_ram_mem3_193_24,
         p_wishbone_bd_ram_mem3_193_25, p_wishbone_bd_ram_mem3_193_26,
         p_wishbone_bd_ram_mem3_193_27, p_wishbone_bd_ram_mem3_193_28,
         p_wishbone_bd_ram_mem3_193_29, p_wishbone_bd_ram_mem3_193_30,
         p_wishbone_bd_ram_mem3_193_31, p_wishbone_bd_ram_mem3_194_24,
         p_wishbone_bd_ram_mem3_194_25, p_wishbone_bd_ram_mem3_194_26,
         p_wishbone_bd_ram_mem3_194_27, p_wishbone_bd_ram_mem3_194_28,
         p_wishbone_bd_ram_mem3_194_29, p_wishbone_bd_ram_mem3_194_30,
         p_wishbone_bd_ram_mem3_194_31, p_wishbone_bd_ram_mem3_195_24,
         p_wishbone_bd_ram_mem3_195_25, p_wishbone_bd_ram_mem3_195_26,
         p_wishbone_bd_ram_mem3_195_27, p_wishbone_bd_ram_mem3_195_28,
         p_wishbone_bd_ram_mem3_195_29, p_wishbone_bd_ram_mem3_195_30,
         p_wishbone_bd_ram_mem3_195_31, p_wishbone_bd_ram_mem3_196_24,
         p_wishbone_bd_ram_mem3_196_25, p_wishbone_bd_ram_mem3_196_26,
         p_wishbone_bd_ram_mem3_196_27, p_wishbone_bd_ram_mem3_196_28,
         p_wishbone_bd_ram_mem3_196_29, p_wishbone_bd_ram_mem3_196_30,
         p_wishbone_bd_ram_mem3_196_31, p_wishbone_bd_ram_mem3_197_24,
         p_wishbone_bd_ram_mem3_197_25, p_wishbone_bd_ram_mem3_197_26,
         p_wishbone_bd_ram_mem3_197_27, p_wishbone_bd_ram_mem3_197_28,
         p_wishbone_bd_ram_mem3_197_29, p_wishbone_bd_ram_mem3_197_30,
         p_wishbone_bd_ram_mem3_197_31, p_wishbone_bd_ram_mem3_198_24,
         p_wishbone_bd_ram_mem3_198_25, p_wishbone_bd_ram_mem3_198_26,
         p_wishbone_bd_ram_mem3_198_27, p_wishbone_bd_ram_mem3_198_28,
         p_wishbone_bd_ram_mem3_198_29, p_wishbone_bd_ram_mem3_198_30,
         p_wishbone_bd_ram_mem3_198_31, p_wishbone_bd_ram_mem3_199_24,
         p_wishbone_bd_ram_mem3_199_25, p_wishbone_bd_ram_mem3_199_26,
         p_wishbone_bd_ram_mem3_199_27, p_wishbone_bd_ram_mem3_199_28,
         p_wishbone_bd_ram_mem3_199_29, p_wishbone_bd_ram_mem3_199_30,
         p_wishbone_bd_ram_mem3_199_31, p_wishbone_bd_ram_mem3_200_24,
         p_wishbone_bd_ram_mem3_200_25, p_wishbone_bd_ram_mem3_200_26,
         p_wishbone_bd_ram_mem3_200_27, p_wishbone_bd_ram_mem3_200_28,
         p_wishbone_bd_ram_mem3_200_29, p_wishbone_bd_ram_mem3_200_30,
         p_wishbone_bd_ram_mem3_200_31, p_wishbone_bd_ram_mem3_201_24,
         p_wishbone_bd_ram_mem3_201_25, p_wishbone_bd_ram_mem3_201_26,
         p_wishbone_bd_ram_mem3_201_27, p_wishbone_bd_ram_mem3_201_28,
         p_wishbone_bd_ram_mem3_201_29, p_wishbone_bd_ram_mem3_201_30,
         p_wishbone_bd_ram_mem3_201_31, p_wishbone_bd_ram_mem3_202_24,
         p_wishbone_bd_ram_mem3_202_25, p_wishbone_bd_ram_mem3_202_26,
         p_wishbone_bd_ram_mem3_202_27, p_wishbone_bd_ram_mem3_202_28,
         p_wishbone_bd_ram_mem3_202_29, p_wishbone_bd_ram_mem3_202_30,
         p_wishbone_bd_ram_mem3_202_31, p_wishbone_bd_ram_mem3_203_24,
         p_wishbone_bd_ram_mem3_203_25, p_wishbone_bd_ram_mem3_203_26,
         p_wishbone_bd_ram_mem3_203_27, p_wishbone_bd_ram_mem3_203_28,
         p_wishbone_bd_ram_mem3_203_29, p_wishbone_bd_ram_mem3_203_30,
         p_wishbone_bd_ram_mem3_203_31, p_wishbone_bd_ram_mem3_204_24,
         p_wishbone_bd_ram_mem3_204_25, p_wishbone_bd_ram_mem3_204_26,
         p_wishbone_bd_ram_mem3_204_27, p_wishbone_bd_ram_mem3_204_28,
         p_wishbone_bd_ram_mem3_204_29, p_wishbone_bd_ram_mem3_204_30,
         p_wishbone_bd_ram_mem3_204_31, p_wishbone_bd_ram_mem3_205_24,
         p_wishbone_bd_ram_mem3_205_25, p_wishbone_bd_ram_mem3_205_26,
         p_wishbone_bd_ram_mem3_205_27, p_wishbone_bd_ram_mem3_205_28,
         p_wishbone_bd_ram_mem3_205_29, p_wishbone_bd_ram_mem3_205_30,
         p_wishbone_bd_ram_mem3_205_31, p_wishbone_bd_ram_mem3_206_24,
         p_wishbone_bd_ram_mem3_206_25, p_wishbone_bd_ram_mem3_206_26,
         p_wishbone_bd_ram_mem3_206_27, p_wishbone_bd_ram_mem3_206_28,
         p_wishbone_bd_ram_mem3_206_29, p_wishbone_bd_ram_mem3_206_30,
         p_wishbone_bd_ram_mem3_206_31, p_wishbone_bd_ram_mem3_207_24,
         p_wishbone_bd_ram_mem3_207_25, p_wishbone_bd_ram_mem3_207_26,
         p_wishbone_bd_ram_mem3_207_27, p_wishbone_bd_ram_mem3_207_28,
         p_wishbone_bd_ram_mem3_207_29, p_wishbone_bd_ram_mem3_207_30,
         p_wishbone_bd_ram_mem3_207_31, p_wishbone_bd_ram_mem3_208_24,
         p_wishbone_bd_ram_mem3_208_25, p_wishbone_bd_ram_mem3_208_26,
         p_wishbone_bd_ram_mem3_208_27, p_wishbone_bd_ram_mem3_208_28,
         p_wishbone_bd_ram_mem3_208_29, p_wishbone_bd_ram_mem3_208_30,
         p_wishbone_bd_ram_mem3_208_31, p_wishbone_bd_ram_mem3_209_24,
         p_wishbone_bd_ram_mem3_209_25, p_wishbone_bd_ram_mem3_209_26,
         p_wishbone_bd_ram_mem3_209_27, p_wishbone_bd_ram_mem3_209_28,
         p_wishbone_bd_ram_mem3_209_29, p_wishbone_bd_ram_mem3_209_30,
         p_wishbone_bd_ram_mem3_209_31, p_wishbone_bd_ram_mem3_210_24,
         p_wishbone_bd_ram_mem3_210_25, p_wishbone_bd_ram_mem3_210_26,
         p_wishbone_bd_ram_mem3_210_27, p_wishbone_bd_ram_mem3_210_28,
         p_wishbone_bd_ram_mem3_210_29, p_wishbone_bd_ram_mem3_210_30,
         p_wishbone_bd_ram_mem3_210_31, p_wishbone_bd_ram_mem3_211_24,
         p_wishbone_bd_ram_mem3_211_25, p_wishbone_bd_ram_mem3_211_26,
         p_wishbone_bd_ram_mem3_211_27, p_wishbone_bd_ram_mem3_211_28,
         p_wishbone_bd_ram_mem3_211_29, p_wishbone_bd_ram_mem3_211_30,
         p_wishbone_bd_ram_mem3_211_31, p_wishbone_bd_ram_mem3_212_24,
         p_wishbone_bd_ram_mem3_212_25, p_wishbone_bd_ram_mem3_212_26,
         p_wishbone_bd_ram_mem3_212_27, p_wishbone_bd_ram_mem3_212_28,
         p_wishbone_bd_ram_mem3_212_29, p_wishbone_bd_ram_mem3_212_30,
         p_wishbone_bd_ram_mem3_212_31, p_wishbone_bd_ram_mem3_213_24,
         p_wishbone_bd_ram_mem3_213_25, p_wishbone_bd_ram_mem3_213_26,
         p_wishbone_bd_ram_mem3_213_27, p_wishbone_bd_ram_mem3_213_28,
         p_wishbone_bd_ram_mem3_213_29, p_wishbone_bd_ram_mem3_213_30,
         p_wishbone_bd_ram_mem3_213_31, p_wishbone_bd_ram_mem3_214_24,
         p_wishbone_bd_ram_mem3_214_25, p_wishbone_bd_ram_mem3_214_26,
         p_wishbone_bd_ram_mem3_214_27, p_wishbone_bd_ram_mem3_214_28,
         p_wishbone_bd_ram_mem3_214_29, p_wishbone_bd_ram_mem3_214_30,
         p_wishbone_bd_ram_mem3_214_31, p_wishbone_bd_ram_mem3_215_24,
         p_wishbone_bd_ram_mem3_215_25, p_wishbone_bd_ram_mem3_215_26,
         p_wishbone_bd_ram_mem3_215_27, p_wishbone_bd_ram_mem3_215_28,
         p_wishbone_bd_ram_mem3_215_29, p_wishbone_bd_ram_mem3_215_30,
         p_wishbone_bd_ram_mem3_215_31, p_wishbone_bd_ram_mem3_216_24,
         p_wishbone_bd_ram_mem3_216_25, p_wishbone_bd_ram_mem3_216_26,
         p_wishbone_bd_ram_mem3_216_27, p_wishbone_bd_ram_mem3_216_28,
         p_wishbone_bd_ram_mem3_216_29, p_wishbone_bd_ram_mem3_216_30,
         p_wishbone_bd_ram_mem3_216_31, p_wishbone_bd_ram_mem3_217_24,
         p_wishbone_bd_ram_mem3_217_25, p_wishbone_bd_ram_mem3_217_26,
         p_wishbone_bd_ram_mem3_217_27, p_wishbone_bd_ram_mem3_217_28,
         p_wishbone_bd_ram_mem3_217_29, p_wishbone_bd_ram_mem3_217_30,
         p_wishbone_bd_ram_mem3_217_31, p_wishbone_bd_ram_mem3_218_24,
         p_wishbone_bd_ram_mem3_218_25, p_wishbone_bd_ram_mem3_218_26,
         p_wishbone_bd_ram_mem3_218_27, p_wishbone_bd_ram_mem3_218_28,
         p_wishbone_bd_ram_mem3_218_29, p_wishbone_bd_ram_mem3_218_30,
         p_wishbone_bd_ram_mem3_218_31, p_wishbone_bd_ram_mem3_219_24,
         p_wishbone_bd_ram_mem3_219_25, p_wishbone_bd_ram_mem3_219_26,
         p_wishbone_bd_ram_mem3_219_27, p_wishbone_bd_ram_mem3_219_28,
         p_wishbone_bd_ram_mem3_219_29, p_wishbone_bd_ram_mem3_219_30,
         p_wishbone_bd_ram_mem3_219_31, p_wishbone_bd_ram_mem3_220_24,
         p_wishbone_bd_ram_mem3_220_25, p_wishbone_bd_ram_mem3_220_26,
         p_wishbone_bd_ram_mem3_220_27, p_wishbone_bd_ram_mem3_220_28,
         p_wishbone_bd_ram_mem3_220_29, p_wishbone_bd_ram_mem3_220_30,
         p_wishbone_bd_ram_mem3_220_31, p_wishbone_bd_ram_mem3_221_24,
         p_wishbone_bd_ram_mem3_221_25, p_wishbone_bd_ram_mem3_221_26,
         p_wishbone_bd_ram_mem3_221_27, p_wishbone_bd_ram_mem3_221_28,
         p_wishbone_bd_ram_mem3_221_29, p_wishbone_bd_ram_mem3_221_30,
         p_wishbone_bd_ram_mem3_221_31, p_wishbone_bd_ram_mem3_222_24,
         p_wishbone_bd_ram_mem3_222_25, p_wishbone_bd_ram_mem3_222_26,
         p_wishbone_bd_ram_mem3_222_27, p_wishbone_bd_ram_mem3_222_28,
         p_wishbone_bd_ram_mem3_222_29, p_wishbone_bd_ram_mem3_222_30,
         p_wishbone_bd_ram_mem3_222_31, p_wishbone_bd_ram_mem3_223_24,
         p_wishbone_bd_ram_mem3_223_25, p_wishbone_bd_ram_mem3_223_26,
         p_wishbone_bd_ram_mem3_223_27, p_wishbone_bd_ram_mem3_223_28,
         p_wishbone_bd_ram_mem3_223_29, p_wishbone_bd_ram_mem3_223_30,
         p_wishbone_bd_ram_mem3_223_31, p_wishbone_bd_ram_mem3_224_24,
         p_wishbone_bd_ram_mem3_224_25, p_wishbone_bd_ram_mem3_224_26,
         p_wishbone_bd_ram_mem3_224_27, p_wishbone_bd_ram_mem3_224_28,
         p_wishbone_bd_ram_mem3_224_29, p_wishbone_bd_ram_mem3_224_30,
         p_wishbone_bd_ram_mem3_224_31, p_wishbone_bd_ram_mem3_225_24,
         p_wishbone_bd_ram_mem3_225_25, p_wishbone_bd_ram_mem3_225_26,
         p_wishbone_bd_ram_mem3_225_27, p_wishbone_bd_ram_mem3_225_28,
         p_wishbone_bd_ram_mem3_225_29, p_wishbone_bd_ram_mem3_225_30,
         p_wishbone_bd_ram_mem3_225_31, p_wishbone_bd_ram_mem3_226_24,
         p_wishbone_bd_ram_mem3_226_25, p_wishbone_bd_ram_mem3_226_26,
         p_wishbone_bd_ram_mem3_226_27, p_wishbone_bd_ram_mem3_226_28,
         p_wishbone_bd_ram_mem3_226_29, p_wishbone_bd_ram_mem3_226_30,
         p_wishbone_bd_ram_mem3_226_31, p_wishbone_bd_ram_mem3_227_24,
         p_wishbone_bd_ram_mem3_227_25, p_wishbone_bd_ram_mem3_227_26,
         p_wishbone_bd_ram_mem3_227_27, p_wishbone_bd_ram_mem3_227_28,
         p_wishbone_bd_ram_mem3_227_29, p_wishbone_bd_ram_mem3_227_30,
         p_wishbone_bd_ram_mem3_227_31, p_wishbone_bd_ram_mem3_228_24,
         p_wishbone_bd_ram_mem3_228_25, p_wishbone_bd_ram_mem3_228_26,
         p_wishbone_bd_ram_mem3_228_27, p_wishbone_bd_ram_mem3_228_28,
         p_wishbone_bd_ram_mem3_228_29, p_wishbone_bd_ram_mem3_228_30,
         p_wishbone_bd_ram_mem3_228_31, p_wishbone_bd_ram_mem3_229_24,
         p_wishbone_bd_ram_mem3_229_25, p_wishbone_bd_ram_mem3_229_26,
         p_wishbone_bd_ram_mem3_229_27, p_wishbone_bd_ram_mem3_229_28,
         p_wishbone_bd_ram_mem3_229_29, p_wishbone_bd_ram_mem3_229_30,
         p_wishbone_bd_ram_mem3_229_31, p_wishbone_bd_ram_mem3_230_24,
         p_wishbone_bd_ram_mem3_230_25, p_wishbone_bd_ram_mem3_230_26,
         p_wishbone_bd_ram_mem3_230_27, p_wishbone_bd_ram_mem3_230_28,
         p_wishbone_bd_ram_mem3_230_29, p_wishbone_bd_ram_mem3_230_30,
         p_wishbone_bd_ram_mem3_230_31, p_wishbone_bd_ram_mem3_231_24,
         p_wishbone_bd_ram_mem3_231_25, p_wishbone_bd_ram_mem3_231_26,
         p_wishbone_bd_ram_mem3_231_27, p_wishbone_bd_ram_mem3_231_28,
         p_wishbone_bd_ram_mem3_231_29, p_wishbone_bd_ram_mem3_231_30,
         p_wishbone_bd_ram_mem3_231_31, p_wishbone_bd_ram_mem3_232_24,
         p_wishbone_bd_ram_mem3_232_25, p_wishbone_bd_ram_mem3_232_26,
         p_wishbone_bd_ram_mem3_232_27, p_wishbone_bd_ram_mem3_232_28,
         p_wishbone_bd_ram_mem3_232_29, p_wishbone_bd_ram_mem3_232_30,
         p_wishbone_bd_ram_mem3_232_31, p_wishbone_bd_ram_mem3_233_24,
         p_wishbone_bd_ram_mem3_233_25, p_wishbone_bd_ram_mem3_233_26,
         p_wishbone_bd_ram_mem3_233_27, p_wishbone_bd_ram_mem3_233_28,
         p_wishbone_bd_ram_mem3_233_29, p_wishbone_bd_ram_mem3_233_30,
         p_wishbone_bd_ram_mem3_233_31, p_wishbone_bd_ram_mem3_234_24,
         p_wishbone_bd_ram_mem3_234_25, p_wishbone_bd_ram_mem3_234_26,
         p_wishbone_bd_ram_mem3_234_27, p_wishbone_bd_ram_mem3_234_28,
         p_wishbone_bd_ram_mem3_234_29, p_wishbone_bd_ram_mem3_234_30,
         p_wishbone_bd_ram_mem3_234_31, p_wishbone_bd_ram_mem3_235_24,
         p_wishbone_bd_ram_mem3_235_25, p_wishbone_bd_ram_mem3_235_26,
         p_wishbone_bd_ram_mem3_235_27, p_wishbone_bd_ram_mem3_235_28,
         p_wishbone_bd_ram_mem3_235_29, p_wishbone_bd_ram_mem3_235_30,
         p_wishbone_bd_ram_mem3_235_31, p_wishbone_bd_ram_mem3_236_24,
         p_wishbone_bd_ram_mem3_236_25, p_wishbone_bd_ram_mem3_236_26,
         p_wishbone_bd_ram_mem3_236_27, p_wishbone_bd_ram_mem3_236_28,
         p_wishbone_bd_ram_mem3_236_29, p_wishbone_bd_ram_mem3_236_30,
         p_wishbone_bd_ram_mem3_236_31, p_wishbone_bd_ram_mem3_237_24,
         p_wishbone_bd_ram_mem3_237_25, p_wishbone_bd_ram_mem3_237_26,
         p_wishbone_bd_ram_mem3_237_27, p_wishbone_bd_ram_mem3_237_28,
         p_wishbone_bd_ram_mem3_237_29, p_wishbone_bd_ram_mem3_237_30,
         p_wishbone_bd_ram_mem3_237_31, p_wishbone_bd_ram_mem3_238_24,
         p_wishbone_bd_ram_mem3_238_25, p_wishbone_bd_ram_mem3_238_26,
         p_wishbone_bd_ram_mem3_238_27, p_wishbone_bd_ram_mem3_238_28,
         p_wishbone_bd_ram_mem3_238_29, p_wishbone_bd_ram_mem3_238_30,
         p_wishbone_bd_ram_mem3_238_31, p_wishbone_bd_ram_mem3_239_24,
         p_wishbone_bd_ram_mem3_239_25, p_wishbone_bd_ram_mem3_239_26,
         p_wishbone_bd_ram_mem3_239_27, p_wishbone_bd_ram_mem3_239_28,
         p_wishbone_bd_ram_mem3_239_29, p_wishbone_bd_ram_mem3_239_30,
         p_wishbone_bd_ram_mem3_239_31, p_wishbone_bd_ram_mem3_240_24,
         p_wishbone_bd_ram_mem3_240_25, p_wishbone_bd_ram_mem3_240_26,
         p_wishbone_bd_ram_mem3_240_27, p_wishbone_bd_ram_mem3_240_28,
         p_wishbone_bd_ram_mem3_240_29, p_wishbone_bd_ram_mem3_240_30,
         p_wishbone_bd_ram_mem3_240_31, p_wishbone_bd_ram_mem3_241_24,
         p_wishbone_bd_ram_mem3_241_25, p_wishbone_bd_ram_mem3_241_26,
         p_wishbone_bd_ram_mem3_241_27, p_wishbone_bd_ram_mem3_241_28,
         p_wishbone_bd_ram_mem3_241_29, p_wishbone_bd_ram_mem3_241_30,
         p_wishbone_bd_ram_mem3_241_31, p_wishbone_bd_ram_mem3_242_24,
         p_wishbone_bd_ram_mem3_242_25, p_wishbone_bd_ram_mem3_242_26,
         p_wishbone_bd_ram_mem3_242_27, p_wishbone_bd_ram_mem3_242_28,
         p_wishbone_bd_ram_mem3_242_29, p_wishbone_bd_ram_mem3_242_30,
         p_wishbone_bd_ram_mem3_242_31, p_wishbone_bd_ram_mem3_243_24,
         p_wishbone_bd_ram_mem3_243_25, p_wishbone_bd_ram_mem3_243_26,
         p_wishbone_bd_ram_mem3_243_27, p_wishbone_bd_ram_mem3_243_28,
         p_wishbone_bd_ram_mem3_243_29, p_wishbone_bd_ram_mem3_243_30,
         p_wishbone_bd_ram_mem3_243_31, p_wishbone_bd_ram_mem3_244_24,
         p_wishbone_bd_ram_mem3_244_25, p_wishbone_bd_ram_mem3_244_26,
         p_wishbone_bd_ram_mem3_244_27, p_wishbone_bd_ram_mem3_244_28,
         p_wishbone_bd_ram_mem3_244_29, p_wishbone_bd_ram_mem3_244_30,
         p_wishbone_bd_ram_mem3_244_31, p_wishbone_bd_ram_mem3_245_24,
         p_wishbone_bd_ram_mem3_245_25, p_wishbone_bd_ram_mem3_245_26,
         p_wishbone_bd_ram_mem3_245_27, p_wishbone_bd_ram_mem3_245_28,
         p_wishbone_bd_ram_mem3_245_29, p_wishbone_bd_ram_mem3_245_30,
         p_wishbone_bd_ram_mem3_245_31, p_wishbone_bd_ram_mem3_246_24,
         p_wishbone_bd_ram_mem3_246_25, p_wishbone_bd_ram_mem3_246_26,
         p_wishbone_bd_ram_mem3_246_27, p_wishbone_bd_ram_mem3_246_28,
         p_wishbone_bd_ram_mem3_246_29, p_wishbone_bd_ram_mem3_246_30,
         p_wishbone_bd_ram_mem3_246_31, p_wishbone_bd_ram_mem3_247_24,
         p_wishbone_bd_ram_mem3_247_25, p_wishbone_bd_ram_mem3_247_26,
         p_wishbone_bd_ram_mem3_247_27, p_wishbone_bd_ram_mem3_247_28,
         p_wishbone_bd_ram_mem3_247_29, p_wishbone_bd_ram_mem3_247_30,
         p_wishbone_bd_ram_mem3_247_31, p_wishbone_bd_ram_mem3_248_24,
         p_wishbone_bd_ram_mem3_248_25, p_wishbone_bd_ram_mem3_248_26,
         p_wishbone_bd_ram_mem3_248_27, p_wishbone_bd_ram_mem3_248_28,
         p_wishbone_bd_ram_mem3_248_29, p_wishbone_bd_ram_mem3_248_30,
         p_wishbone_bd_ram_mem3_248_31, p_wishbone_bd_ram_mem3_249_24,
         p_wishbone_bd_ram_mem3_249_25, p_wishbone_bd_ram_mem3_249_26,
         p_wishbone_bd_ram_mem3_249_27, p_wishbone_bd_ram_mem3_249_28,
         p_wishbone_bd_ram_mem3_249_29, p_wishbone_bd_ram_mem3_249_30,
         p_wishbone_bd_ram_mem3_249_31, p_wishbone_bd_ram_mem3_250_24,
         p_wishbone_bd_ram_mem3_250_25, p_wishbone_bd_ram_mem3_250_26,
         p_wishbone_bd_ram_mem3_250_27, p_wishbone_bd_ram_mem3_250_28,
         p_wishbone_bd_ram_mem3_250_29, p_wishbone_bd_ram_mem3_250_30,
         p_wishbone_bd_ram_mem3_250_31, p_wishbone_bd_ram_mem3_251_24,
         p_wishbone_bd_ram_mem3_251_25, p_wishbone_bd_ram_mem3_251_26,
         p_wishbone_bd_ram_mem3_251_27, p_wishbone_bd_ram_mem3_251_28,
         p_wishbone_bd_ram_mem3_251_29, p_wishbone_bd_ram_mem3_251_30,
         p_wishbone_bd_ram_mem3_251_31, p_wishbone_bd_ram_mem3_252_24,
         p_wishbone_bd_ram_mem3_252_25, p_wishbone_bd_ram_mem3_252_26,
         p_wishbone_bd_ram_mem3_252_27, p_wishbone_bd_ram_mem3_252_28,
         p_wishbone_bd_ram_mem3_252_29, p_wishbone_bd_ram_mem3_252_30,
         p_wishbone_bd_ram_mem3_252_31, p_wishbone_bd_ram_mem3_253_24,
         p_wishbone_bd_ram_mem3_253_25, p_wishbone_bd_ram_mem3_253_26,
         p_wishbone_bd_ram_mem3_253_27, p_wishbone_bd_ram_mem3_253_28,
         p_wishbone_bd_ram_mem3_253_29, p_wishbone_bd_ram_mem3_253_30,
         p_wishbone_bd_ram_mem3_253_31, p_wishbone_bd_ram_mem3_254_24,
         p_wishbone_bd_ram_mem3_254_25, p_wishbone_bd_ram_mem3_254_26,
         p_wishbone_bd_ram_mem3_254_27, p_wishbone_bd_ram_mem3_254_28,
         p_wishbone_bd_ram_mem3_254_29, p_wishbone_bd_ram_mem3_254_30,
         p_wishbone_bd_ram_mem3_254_31, p_wishbone_bd_ram_mem3_255_24,
         p_wishbone_bd_ram_mem3_255_25, p_wishbone_bd_ram_mem3_255_26,
         p_wishbone_bd_ram_mem3_255_27, p_wishbone_bd_ram_mem3_255_28,
         p_wishbone_bd_ram_mem3_255_29, p_wishbone_bd_ram_mem3_255_30,
         p_wishbone_bd_ram_mem3_255_31, p_wishbone_bd_ram_mem1_0_8,
         p_wishbone_bd_ram_mem1_0_9, p_wishbone_bd_ram_mem1_0_10,
         p_wishbone_bd_ram_mem1_0_11, p_wishbone_bd_ram_mem1_0_12,
         p_wishbone_bd_ram_mem1_0_13, p_wishbone_bd_ram_mem1_0_14,
         p_wishbone_bd_ram_mem1_0_15, p_wishbone_bd_ram_mem1_1_8,
         p_wishbone_bd_ram_mem1_1_9, p_wishbone_bd_ram_mem1_1_10,
         p_wishbone_bd_ram_mem1_1_11, p_wishbone_bd_ram_mem1_1_12,
         p_wishbone_bd_ram_mem1_1_13, p_wishbone_bd_ram_mem1_1_14,
         p_wishbone_bd_ram_mem1_1_15, p_wishbone_bd_ram_mem1_2_8,
         p_wishbone_bd_ram_mem1_2_9, p_wishbone_bd_ram_mem1_2_10,
         p_wishbone_bd_ram_mem1_2_11, p_wishbone_bd_ram_mem1_2_12,
         p_wishbone_bd_ram_mem1_2_13, p_wishbone_bd_ram_mem1_2_14,
         p_wishbone_bd_ram_mem1_2_15, p_wishbone_bd_ram_mem1_3_8,
         p_wishbone_bd_ram_mem1_3_9, p_wishbone_bd_ram_mem1_3_10,
         p_wishbone_bd_ram_mem1_3_11, p_wishbone_bd_ram_mem1_3_12,
         p_wishbone_bd_ram_mem1_3_13, p_wishbone_bd_ram_mem1_3_14,
         p_wishbone_bd_ram_mem1_3_15, p_wishbone_bd_ram_mem1_4_8,
         p_wishbone_bd_ram_mem1_4_9, p_wishbone_bd_ram_mem1_4_10,
         p_wishbone_bd_ram_mem1_4_11, p_wishbone_bd_ram_mem1_4_12,
         p_wishbone_bd_ram_mem1_4_13, p_wishbone_bd_ram_mem1_4_14,
         p_wishbone_bd_ram_mem1_4_15, p_wishbone_bd_ram_mem1_5_8,
         p_wishbone_bd_ram_mem1_5_9, p_wishbone_bd_ram_mem1_5_10,
         p_wishbone_bd_ram_mem1_5_11, p_wishbone_bd_ram_mem1_5_12,
         p_wishbone_bd_ram_mem1_5_13, p_wishbone_bd_ram_mem1_5_14,
         p_wishbone_bd_ram_mem1_5_15, p_wishbone_bd_ram_mem1_6_8,
         p_wishbone_bd_ram_mem1_6_9, p_wishbone_bd_ram_mem1_6_10,
         p_wishbone_bd_ram_mem1_6_11, p_wishbone_bd_ram_mem1_6_12,
         p_wishbone_bd_ram_mem1_6_13, p_wishbone_bd_ram_mem1_6_14,
         p_wishbone_bd_ram_mem1_6_15, p_wishbone_bd_ram_mem1_7_8,
         p_wishbone_bd_ram_mem1_7_9, p_wishbone_bd_ram_mem1_7_10,
         p_wishbone_bd_ram_mem1_7_11, p_wishbone_bd_ram_mem1_7_12,
         p_wishbone_bd_ram_mem1_7_13, p_wishbone_bd_ram_mem1_7_14,
         p_wishbone_bd_ram_mem1_7_15, p_wishbone_bd_ram_mem1_8_8,
         p_wishbone_bd_ram_mem1_8_9, p_wishbone_bd_ram_mem1_8_10,
         p_wishbone_bd_ram_mem1_8_11, p_wishbone_bd_ram_mem1_8_12,
         p_wishbone_bd_ram_mem1_8_13, p_wishbone_bd_ram_mem1_8_14,
         p_wishbone_bd_ram_mem1_8_15, p_wishbone_bd_ram_mem1_9_8,
         p_wishbone_bd_ram_mem1_9_9, p_wishbone_bd_ram_mem1_9_10,
         p_wishbone_bd_ram_mem1_9_11, p_wishbone_bd_ram_mem1_9_12,
         p_wishbone_bd_ram_mem1_9_13, p_wishbone_bd_ram_mem1_9_14,
         p_wishbone_bd_ram_mem1_9_15, p_wishbone_bd_ram_mem1_10_8,
         p_wishbone_bd_ram_mem1_10_9, p_wishbone_bd_ram_mem1_10_10,
         p_wishbone_bd_ram_mem1_10_11, p_wishbone_bd_ram_mem1_10_12,
         p_wishbone_bd_ram_mem1_10_13, p_wishbone_bd_ram_mem1_10_14,
         p_wishbone_bd_ram_mem1_10_15, p_wishbone_bd_ram_mem1_11_8,
         p_wishbone_bd_ram_mem1_11_9, p_wishbone_bd_ram_mem1_11_10,
         p_wishbone_bd_ram_mem1_11_11, p_wishbone_bd_ram_mem1_11_12,
         p_wishbone_bd_ram_mem1_11_13, p_wishbone_bd_ram_mem1_11_14,
         p_wishbone_bd_ram_mem1_11_15, p_wishbone_bd_ram_mem1_12_8,
         p_wishbone_bd_ram_mem1_12_9, p_wishbone_bd_ram_mem1_12_10,
         p_wishbone_bd_ram_mem1_12_11, p_wishbone_bd_ram_mem1_12_12,
         p_wishbone_bd_ram_mem1_12_13, p_wishbone_bd_ram_mem1_12_14,
         p_wishbone_bd_ram_mem1_12_15, p_wishbone_bd_ram_mem1_13_8,
         p_wishbone_bd_ram_mem1_13_9, p_wishbone_bd_ram_mem1_13_10,
         p_wishbone_bd_ram_mem1_13_11, p_wishbone_bd_ram_mem1_13_12,
         p_wishbone_bd_ram_mem1_13_13, p_wishbone_bd_ram_mem1_13_14,
         p_wishbone_bd_ram_mem1_13_15, p_wishbone_bd_ram_mem1_14_8,
         p_wishbone_bd_ram_mem1_14_9, p_wishbone_bd_ram_mem1_14_10,
         p_wishbone_bd_ram_mem1_14_11, p_wishbone_bd_ram_mem1_14_12,
         p_wishbone_bd_ram_mem1_14_13, p_wishbone_bd_ram_mem1_14_14,
         p_wishbone_bd_ram_mem1_14_15, p_wishbone_bd_ram_mem1_15_8,
         p_wishbone_bd_ram_mem1_15_9, p_wishbone_bd_ram_mem1_15_10,
         p_wishbone_bd_ram_mem1_15_11, p_wishbone_bd_ram_mem1_15_12,
         p_wishbone_bd_ram_mem1_15_13, p_wishbone_bd_ram_mem1_15_14,
         p_wishbone_bd_ram_mem1_15_15, p_wishbone_bd_ram_mem1_16_8,
         p_wishbone_bd_ram_mem1_16_9, p_wishbone_bd_ram_mem1_16_10,
         p_wishbone_bd_ram_mem1_16_11, p_wishbone_bd_ram_mem1_16_12,
         p_wishbone_bd_ram_mem1_16_13, p_wishbone_bd_ram_mem1_16_14,
         p_wishbone_bd_ram_mem1_16_15, p_wishbone_bd_ram_mem1_17_8,
         p_wishbone_bd_ram_mem1_17_9, p_wishbone_bd_ram_mem1_17_10,
         p_wishbone_bd_ram_mem1_17_11, p_wishbone_bd_ram_mem1_17_12,
         p_wishbone_bd_ram_mem1_17_13, p_wishbone_bd_ram_mem1_17_14,
         p_wishbone_bd_ram_mem1_17_15, p_wishbone_bd_ram_mem1_18_8,
         p_wishbone_bd_ram_mem1_18_9, p_wishbone_bd_ram_mem1_18_10,
         p_wishbone_bd_ram_mem1_18_11, p_wishbone_bd_ram_mem1_18_12,
         p_wishbone_bd_ram_mem1_18_13, p_wishbone_bd_ram_mem1_18_14,
         p_wishbone_bd_ram_mem1_18_15, p_wishbone_bd_ram_mem1_19_8,
         p_wishbone_bd_ram_mem1_19_9, p_wishbone_bd_ram_mem1_19_10,
         p_wishbone_bd_ram_mem1_19_11, p_wishbone_bd_ram_mem1_19_12,
         p_wishbone_bd_ram_mem1_19_13, p_wishbone_bd_ram_mem1_19_14,
         p_wishbone_bd_ram_mem1_19_15, p_wishbone_bd_ram_mem1_20_8,
         p_wishbone_bd_ram_mem1_20_9, p_wishbone_bd_ram_mem1_20_10,
         p_wishbone_bd_ram_mem1_20_11, p_wishbone_bd_ram_mem1_20_12,
         p_wishbone_bd_ram_mem1_20_13, p_wishbone_bd_ram_mem1_20_14,
         p_wishbone_bd_ram_mem1_20_15, p_wishbone_bd_ram_mem1_21_8,
         p_wishbone_bd_ram_mem1_21_9, p_wishbone_bd_ram_mem1_21_10,
         p_wishbone_bd_ram_mem1_21_11, p_wishbone_bd_ram_mem1_21_12,
         p_wishbone_bd_ram_mem1_21_13, p_wishbone_bd_ram_mem1_21_14,
         p_wishbone_bd_ram_mem1_21_15, p_wishbone_bd_ram_mem1_22_8,
         p_wishbone_bd_ram_mem1_22_9, p_wishbone_bd_ram_mem1_22_10,
         p_wishbone_bd_ram_mem1_22_11, p_wishbone_bd_ram_mem1_22_12,
         p_wishbone_bd_ram_mem1_22_13, p_wishbone_bd_ram_mem1_22_14,
         p_wishbone_bd_ram_mem1_22_15, p_wishbone_bd_ram_mem1_23_8,
         p_wishbone_bd_ram_mem1_23_9, p_wishbone_bd_ram_mem1_23_10,
         p_wishbone_bd_ram_mem1_23_11, p_wishbone_bd_ram_mem1_23_12,
         p_wishbone_bd_ram_mem1_23_13, p_wishbone_bd_ram_mem1_23_14,
         p_wishbone_bd_ram_mem1_23_15, p_wishbone_bd_ram_mem1_24_8,
         p_wishbone_bd_ram_mem1_24_9, p_wishbone_bd_ram_mem1_24_10,
         p_wishbone_bd_ram_mem1_24_11, p_wishbone_bd_ram_mem1_24_12,
         p_wishbone_bd_ram_mem1_24_13, p_wishbone_bd_ram_mem1_24_14,
         p_wishbone_bd_ram_mem1_24_15, p_wishbone_bd_ram_mem1_25_8,
         p_wishbone_bd_ram_mem1_25_9, p_wishbone_bd_ram_mem1_25_10,
         p_wishbone_bd_ram_mem1_25_11, p_wishbone_bd_ram_mem1_25_12,
         p_wishbone_bd_ram_mem1_25_13, p_wishbone_bd_ram_mem1_25_14,
         p_wishbone_bd_ram_mem1_25_15, p_wishbone_bd_ram_mem1_26_8,
         p_wishbone_bd_ram_mem1_26_9, p_wishbone_bd_ram_mem1_26_10,
         p_wishbone_bd_ram_mem1_26_11, p_wishbone_bd_ram_mem1_26_12,
         p_wishbone_bd_ram_mem1_26_13, p_wishbone_bd_ram_mem1_26_14,
         p_wishbone_bd_ram_mem1_26_15, p_wishbone_bd_ram_mem1_27_8,
         p_wishbone_bd_ram_mem1_27_9, p_wishbone_bd_ram_mem1_27_10,
         p_wishbone_bd_ram_mem1_27_11, p_wishbone_bd_ram_mem1_27_12,
         p_wishbone_bd_ram_mem1_27_13, p_wishbone_bd_ram_mem1_27_14,
         p_wishbone_bd_ram_mem1_27_15, p_wishbone_bd_ram_mem1_28_8,
         p_wishbone_bd_ram_mem1_28_9, p_wishbone_bd_ram_mem1_28_10,
         p_wishbone_bd_ram_mem1_28_11, p_wishbone_bd_ram_mem1_28_12,
         p_wishbone_bd_ram_mem1_28_13, p_wishbone_bd_ram_mem1_28_14,
         p_wishbone_bd_ram_mem1_28_15, p_wishbone_bd_ram_mem1_29_8,
         p_wishbone_bd_ram_mem1_29_9, p_wishbone_bd_ram_mem1_29_10,
         p_wishbone_bd_ram_mem1_29_11, p_wishbone_bd_ram_mem1_29_12,
         p_wishbone_bd_ram_mem1_29_13, p_wishbone_bd_ram_mem1_29_14,
         p_wishbone_bd_ram_mem1_29_15, p_wishbone_bd_ram_mem1_30_8,
         p_wishbone_bd_ram_mem1_30_9, p_wishbone_bd_ram_mem1_30_10,
         p_wishbone_bd_ram_mem1_30_11, p_wishbone_bd_ram_mem1_30_12,
         p_wishbone_bd_ram_mem1_30_13, p_wishbone_bd_ram_mem1_30_14,
         p_wishbone_bd_ram_mem1_30_15, p_wishbone_bd_ram_mem1_31_8,
         p_wishbone_bd_ram_mem1_31_9, p_wishbone_bd_ram_mem1_31_10,
         p_wishbone_bd_ram_mem1_31_11, p_wishbone_bd_ram_mem1_31_12,
         p_wishbone_bd_ram_mem1_31_13, p_wishbone_bd_ram_mem1_31_14,
         p_wishbone_bd_ram_mem1_31_15, p_wishbone_bd_ram_mem1_32_8,
         p_wishbone_bd_ram_mem1_32_9, p_wishbone_bd_ram_mem1_32_10,
         p_wishbone_bd_ram_mem1_32_11, p_wishbone_bd_ram_mem1_32_12,
         p_wishbone_bd_ram_mem1_32_13, p_wishbone_bd_ram_mem1_32_14,
         p_wishbone_bd_ram_mem1_32_15, p_wishbone_bd_ram_mem1_33_8,
         p_wishbone_bd_ram_mem1_33_9, p_wishbone_bd_ram_mem1_33_10,
         p_wishbone_bd_ram_mem1_33_11, p_wishbone_bd_ram_mem1_33_12,
         p_wishbone_bd_ram_mem1_33_13, p_wishbone_bd_ram_mem1_33_14,
         p_wishbone_bd_ram_mem1_33_15, p_wishbone_bd_ram_mem1_34_8,
         p_wishbone_bd_ram_mem1_34_9, p_wishbone_bd_ram_mem1_34_10,
         p_wishbone_bd_ram_mem1_34_11, p_wishbone_bd_ram_mem1_34_12,
         p_wishbone_bd_ram_mem1_34_13, p_wishbone_bd_ram_mem1_34_14,
         p_wishbone_bd_ram_mem1_34_15, p_wishbone_bd_ram_mem1_35_8,
         p_wishbone_bd_ram_mem1_35_9, p_wishbone_bd_ram_mem1_35_10,
         p_wishbone_bd_ram_mem1_35_11, p_wishbone_bd_ram_mem1_35_12,
         p_wishbone_bd_ram_mem1_35_13, p_wishbone_bd_ram_mem1_35_14,
         p_wishbone_bd_ram_mem1_35_15, p_wishbone_bd_ram_mem1_36_8,
         p_wishbone_bd_ram_mem1_36_9, p_wishbone_bd_ram_mem1_36_10,
         p_wishbone_bd_ram_mem1_36_11, p_wishbone_bd_ram_mem1_36_12,
         p_wishbone_bd_ram_mem1_36_13, p_wishbone_bd_ram_mem1_36_14,
         p_wishbone_bd_ram_mem1_36_15, p_wishbone_bd_ram_mem1_37_8,
         p_wishbone_bd_ram_mem1_37_9, p_wishbone_bd_ram_mem1_37_10,
         p_wishbone_bd_ram_mem1_37_11, p_wishbone_bd_ram_mem1_37_12,
         p_wishbone_bd_ram_mem1_37_13, p_wishbone_bd_ram_mem1_37_14,
         p_wishbone_bd_ram_mem1_37_15, p_wishbone_bd_ram_mem1_38_8,
         p_wishbone_bd_ram_mem1_38_9, p_wishbone_bd_ram_mem1_38_10,
         p_wishbone_bd_ram_mem1_38_11, p_wishbone_bd_ram_mem1_38_12,
         p_wishbone_bd_ram_mem1_38_13, p_wishbone_bd_ram_mem1_38_14,
         p_wishbone_bd_ram_mem1_38_15, p_wishbone_bd_ram_mem1_39_8,
         p_wishbone_bd_ram_mem1_39_9, p_wishbone_bd_ram_mem1_39_10,
         p_wishbone_bd_ram_mem1_39_11, p_wishbone_bd_ram_mem1_39_12,
         p_wishbone_bd_ram_mem1_39_13, p_wishbone_bd_ram_mem1_39_14,
         p_wishbone_bd_ram_mem1_39_15, p_wishbone_bd_ram_mem1_40_8,
         p_wishbone_bd_ram_mem1_40_9, p_wishbone_bd_ram_mem1_40_10,
         p_wishbone_bd_ram_mem1_40_11, p_wishbone_bd_ram_mem1_40_12,
         p_wishbone_bd_ram_mem1_40_13, p_wishbone_bd_ram_mem1_40_14,
         p_wishbone_bd_ram_mem1_40_15, p_wishbone_bd_ram_mem1_41_8,
         p_wishbone_bd_ram_mem1_41_9, p_wishbone_bd_ram_mem1_41_10,
         p_wishbone_bd_ram_mem1_41_11, p_wishbone_bd_ram_mem1_41_12,
         p_wishbone_bd_ram_mem1_41_13, p_wishbone_bd_ram_mem1_41_14,
         p_wishbone_bd_ram_mem1_41_15, p_wishbone_bd_ram_mem1_42_8,
         p_wishbone_bd_ram_mem1_42_9, p_wishbone_bd_ram_mem1_42_10,
         p_wishbone_bd_ram_mem1_42_11, p_wishbone_bd_ram_mem1_42_12,
         p_wishbone_bd_ram_mem1_42_13, p_wishbone_bd_ram_mem1_42_14,
         p_wishbone_bd_ram_mem1_42_15, p_wishbone_bd_ram_mem1_43_8,
         p_wishbone_bd_ram_mem1_43_9, p_wishbone_bd_ram_mem1_43_10,
         p_wishbone_bd_ram_mem1_43_11, p_wishbone_bd_ram_mem1_43_12,
         p_wishbone_bd_ram_mem1_43_13, p_wishbone_bd_ram_mem1_43_14,
         p_wishbone_bd_ram_mem1_43_15, p_wishbone_bd_ram_mem1_44_8,
         p_wishbone_bd_ram_mem1_44_9, p_wishbone_bd_ram_mem1_44_10,
         p_wishbone_bd_ram_mem1_44_11, p_wishbone_bd_ram_mem1_44_12,
         p_wishbone_bd_ram_mem1_44_13, p_wishbone_bd_ram_mem1_44_14,
         p_wishbone_bd_ram_mem1_44_15, p_wishbone_bd_ram_mem1_45_8,
         p_wishbone_bd_ram_mem1_45_9, p_wishbone_bd_ram_mem1_45_10,
         p_wishbone_bd_ram_mem1_45_11, p_wishbone_bd_ram_mem1_45_12,
         p_wishbone_bd_ram_mem1_45_13, p_wishbone_bd_ram_mem1_45_14,
         p_wishbone_bd_ram_mem1_45_15, p_wishbone_bd_ram_mem1_46_8,
         p_wishbone_bd_ram_mem1_46_9, p_wishbone_bd_ram_mem1_46_10,
         p_wishbone_bd_ram_mem1_46_11, p_wishbone_bd_ram_mem1_46_12,
         p_wishbone_bd_ram_mem1_46_13, p_wishbone_bd_ram_mem1_46_14,
         p_wishbone_bd_ram_mem1_46_15, p_wishbone_bd_ram_mem1_47_8,
         p_wishbone_bd_ram_mem1_47_9, p_wishbone_bd_ram_mem1_47_10,
         p_wishbone_bd_ram_mem1_47_11, p_wishbone_bd_ram_mem1_47_12,
         p_wishbone_bd_ram_mem1_47_13, p_wishbone_bd_ram_mem1_47_14,
         p_wishbone_bd_ram_mem1_47_15, p_wishbone_bd_ram_mem1_48_8,
         p_wishbone_bd_ram_mem1_48_9, p_wishbone_bd_ram_mem1_48_10,
         p_wishbone_bd_ram_mem1_48_11, p_wishbone_bd_ram_mem1_48_12,
         p_wishbone_bd_ram_mem1_48_13, p_wishbone_bd_ram_mem1_48_14,
         p_wishbone_bd_ram_mem1_48_15, p_wishbone_bd_ram_mem1_49_8,
         p_wishbone_bd_ram_mem1_49_9, p_wishbone_bd_ram_mem1_49_10,
         p_wishbone_bd_ram_mem1_49_11, p_wishbone_bd_ram_mem1_49_12,
         p_wishbone_bd_ram_mem1_49_13, p_wishbone_bd_ram_mem1_49_14,
         p_wishbone_bd_ram_mem1_49_15, p_wishbone_bd_ram_mem1_50_8,
         p_wishbone_bd_ram_mem1_50_9, p_wishbone_bd_ram_mem1_50_10,
         p_wishbone_bd_ram_mem1_50_11, p_wishbone_bd_ram_mem1_50_12,
         p_wishbone_bd_ram_mem1_50_13, p_wishbone_bd_ram_mem1_50_14,
         p_wishbone_bd_ram_mem1_50_15, p_wishbone_bd_ram_mem1_51_8,
         p_wishbone_bd_ram_mem1_51_9, p_wishbone_bd_ram_mem1_51_10,
         p_wishbone_bd_ram_mem1_51_11, p_wishbone_bd_ram_mem1_51_12,
         p_wishbone_bd_ram_mem1_51_13, p_wishbone_bd_ram_mem1_51_14,
         p_wishbone_bd_ram_mem1_51_15, p_wishbone_bd_ram_mem1_52_8,
         p_wishbone_bd_ram_mem1_52_9, p_wishbone_bd_ram_mem1_52_10,
         p_wishbone_bd_ram_mem1_52_11, p_wishbone_bd_ram_mem1_52_12,
         p_wishbone_bd_ram_mem1_52_13, p_wishbone_bd_ram_mem1_52_14,
         p_wishbone_bd_ram_mem1_52_15, p_wishbone_bd_ram_mem1_53_8,
         p_wishbone_bd_ram_mem1_53_9, p_wishbone_bd_ram_mem1_53_10,
         p_wishbone_bd_ram_mem1_53_11, p_wishbone_bd_ram_mem1_53_12,
         p_wishbone_bd_ram_mem1_53_13, p_wishbone_bd_ram_mem1_53_14,
         p_wishbone_bd_ram_mem1_53_15, p_wishbone_bd_ram_mem1_54_8,
         p_wishbone_bd_ram_mem1_54_9, p_wishbone_bd_ram_mem1_54_10,
         p_wishbone_bd_ram_mem1_54_11, p_wishbone_bd_ram_mem1_54_12,
         p_wishbone_bd_ram_mem1_54_13, p_wishbone_bd_ram_mem1_54_14,
         p_wishbone_bd_ram_mem1_54_15, p_wishbone_bd_ram_mem1_55_8,
         p_wishbone_bd_ram_mem1_55_9, p_wishbone_bd_ram_mem1_55_10,
         p_wishbone_bd_ram_mem1_55_11, p_wishbone_bd_ram_mem1_55_12,
         p_wishbone_bd_ram_mem1_55_13, p_wishbone_bd_ram_mem1_55_14,
         p_wishbone_bd_ram_mem1_55_15, p_wishbone_bd_ram_mem1_56_8,
         p_wishbone_bd_ram_mem1_56_9, p_wishbone_bd_ram_mem1_56_10,
         p_wishbone_bd_ram_mem1_56_11, p_wishbone_bd_ram_mem1_56_12,
         p_wishbone_bd_ram_mem1_56_13, p_wishbone_bd_ram_mem1_56_14,
         p_wishbone_bd_ram_mem1_56_15, p_wishbone_bd_ram_mem1_57_8,
         p_wishbone_bd_ram_mem1_57_9, p_wishbone_bd_ram_mem1_57_10,
         p_wishbone_bd_ram_mem1_57_11, p_wishbone_bd_ram_mem1_57_12,
         p_wishbone_bd_ram_mem1_57_13, p_wishbone_bd_ram_mem1_57_14,
         p_wishbone_bd_ram_mem1_57_15, p_wishbone_bd_ram_mem1_58_8,
         p_wishbone_bd_ram_mem1_58_9, p_wishbone_bd_ram_mem1_58_10,
         p_wishbone_bd_ram_mem1_58_11, p_wishbone_bd_ram_mem1_58_12,
         p_wishbone_bd_ram_mem1_58_13, p_wishbone_bd_ram_mem1_58_14,
         p_wishbone_bd_ram_mem1_58_15, p_wishbone_bd_ram_mem1_59_8,
         p_wishbone_bd_ram_mem1_59_9, p_wishbone_bd_ram_mem1_59_10,
         p_wishbone_bd_ram_mem1_59_11, p_wishbone_bd_ram_mem1_59_12,
         p_wishbone_bd_ram_mem1_59_13, p_wishbone_bd_ram_mem1_59_14,
         p_wishbone_bd_ram_mem1_59_15, p_wishbone_bd_ram_mem1_60_8,
         p_wishbone_bd_ram_mem1_60_9, p_wishbone_bd_ram_mem1_60_10,
         p_wishbone_bd_ram_mem1_60_11, p_wishbone_bd_ram_mem1_60_12,
         p_wishbone_bd_ram_mem1_60_13, p_wishbone_bd_ram_mem1_60_14,
         p_wishbone_bd_ram_mem1_60_15, p_wishbone_bd_ram_mem1_61_8,
         p_wishbone_bd_ram_mem1_61_9, p_wishbone_bd_ram_mem1_61_10,
         p_wishbone_bd_ram_mem1_61_11, p_wishbone_bd_ram_mem1_61_12,
         p_wishbone_bd_ram_mem1_61_13, p_wishbone_bd_ram_mem1_61_14,
         p_wishbone_bd_ram_mem1_61_15, p_wishbone_bd_ram_mem1_62_8,
         p_wishbone_bd_ram_mem1_62_9, p_wishbone_bd_ram_mem1_62_10,
         p_wishbone_bd_ram_mem1_62_11, p_wishbone_bd_ram_mem1_62_12,
         p_wishbone_bd_ram_mem1_62_13, p_wishbone_bd_ram_mem1_62_14,
         p_wishbone_bd_ram_mem1_62_15, p_wishbone_bd_ram_mem1_63_8,
         p_wishbone_bd_ram_mem1_63_9, p_wishbone_bd_ram_mem1_63_10,
         p_wishbone_bd_ram_mem1_63_11, p_wishbone_bd_ram_mem1_63_12,
         p_wishbone_bd_ram_mem1_63_13, p_wishbone_bd_ram_mem1_63_14,
         p_wishbone_bd_ram_mem1_63_15, p_wishbone_bd_ram_mem1_64_8,
         p_wishbone_bd_ram_mem1_64_9, p_wishbone_bd_ram_mem1_64_10,
         p_wishbone_bd_ram_mem1_64_11, p_wishbone_bd_ram_mem1_64_12,
         p_wishbone_bd_ram_mem1_64_13, p_wishbone_bd_ram_mem1_64_14,
         p_wishbone_bd_ram_mem1_64_15, p_wishbone_bd_ram_mem1_65_8,
         p_wishbone_bd_ram_mem1_65_9, p_wishbone_bd_ram_mem1_65_10,
         p_wishbone_bd_ram_mem1_65_11, p_wishbone_bd_ram_mem1_65_12,
         p_wishbone_bd_ram_mem1_65_13, p_wishbone_bd_ram_mem1_65_14,
         p_wishbone_bd_ram_mem1_65_15, p_wishbone_bd_ram_mem1_66_8,
         p_wishbone_bd_ram_mem1_66_9, p_wishbone_bd_ram_mem1_66_10,
         p_wishbone_bd_ram_mem1_66_11, p_wishbone_bd_ram_mem1_66_12,
         p_wishbone_bd_ram_mem1_66_13, p_wishbone_bd_ram_mem1_66_14,
         p_wishbone_bd_ram_mem1_66_15, p_wishbone_bd_ram_mem1_67_8,
         p_wishbone_bd_ram_mem1_67_9, p_wishbone_bd_ram_mem1_67_10,
         p_wishbone_bd_ram_mem1_67_11, p_wishbone_bd_ram_mem1_67_12,
         p_wishbone_bd_ram_mem1_67_13, p_wishbone_bd_ram_mem1_67_14,
         p_wishbone_bd_ram_mem1_67_15, p_wishbone_bd_ram_mem1_68_8,
         p_wishbone_bd_ram_mem1_68_9, p_wishbone_bd_ram_mem1_68_10,
         p_wishbone_bd_ram_mem1_68_11, p_wishbone_bd_ram_mem1_68_12,
         p_wishbone_bd_ram_mem1_68_13, p_wishbone_bd_ram_mem1_68_14,
         p_wishbone_bd_ram_mem1_68_15, p_wishbone_bd_ram_mem1_69_8,
         p_wishbone_bd_ram_mem1_69_9, p_wishbone_bd_ram_mem1_69_10,
         p_wishbone_bd_ram_mem1_69_11, p_wishbone_bd_ram_mem1_69_12,
         p_wishbone_bd_ram_mem1_69_13, p_wishbone_bd_ram_mem1_69_14,
         p_wishbone_bd_ram_mem1_69_15, p_wishbone_bd_ram_mem1_70_8,
         p_wishbone_bd_ram_mem1_70_9, p_wishbone_bd_ram_mem1_70_10,
         p_wishbone_bd_ram_mem1_70_11, p_wishbone_bd_ram_mem1_70_12,
         p_wishbone_bd_ram_mem1_70_13, p_wishbone_bd_ram_mem1_70_14,
         p_wishbone_bd_ram_mem1_70_15, p_wishbone_bd_ram_mem1_71_8,
         p_wishbone_bd_ram_mem1_71_9, p_wishbone_bd_ram_mem1_71_10,
         p_wishbone_bd_ram_mem1_71_11, p_wishbone_bd_ram_mem1_71_12,
         p_wishbone_bd_ram_mem1_71_13, p_wishbone_bd_ram_mem1_71_14,
         p_wishbone_bd_ram_mem1_71_15, p_wishbone_bd_ram_mem1_72_8,
         p_wishbone_bd_ram_mem1_72_9, p_wishbone_bd_ram_mem1_72_10,
         p_wishbone_bd_ram_mem1_72_11, p_wishbone_bd_ram_mem1_72_12,
         p_wishbone_bd_ram_mem1_72_13, p_wishbone_bd_ram_mem1_72_14,
         p_wishbone_bd_ram_mem1_72_15, p_wishbone_bd_ram_mem1_73_8,
         p_wishbone_bd_ram_mem1_73_9, p_wishbone_bd_ram_mem1_73_10,
         p_wishbone_bd_ram_mem1_73_11, p_wishbone_bd_ram_mem1_73_12,
         p_wishbone_bd_ram_mem1_73_13, p_wishbone_bd_ram_mem1_73_14,
         p_wishbone_bd_ram_mem1_73_15, p_wishbone_bd_ram_mem1_74_8,
         p_wishbone_bd_ram_mem1_74_9, p_wishbone_bd_ram_mem1_74_10,
         p_wishbone_bd_ram_mem1_74_11, p_wishbone_bd_ram_mem1_74_12,
         p_wishbone_bd_ram_mem1_74_13, p_wishbone_bd_ram_mem1_74_14,
         p_wishbone_bd_ram_mem1_74_15, p_wishbone_bd_ram_mem1_75_8,
         p_wishbone_bd_ram_mem1_75_9, p_wishbone_bd_ram_mem1_75_10,
         p_wishbone_bd_ram_mem1_75_11, p_wishbone_bd_ram_mem1_75_12,
         p_wishbone_bd_ram_mem1_75_13, p_wishbone_bd_ram_mem1_75_14,
         p_wishbone_bd_ram_mem1_75_15, p_wishbone_bd_ram_mem1_76_8,
         p_wishbone_bd_ram_mem1_76_9, p_wishbone_bd_ram_mem1_76_10,
         p_wishbone_bd_ram_mem1_76_11, p_wishbone_bd_ram_mem1_76_12,
         p_wishbone_bd_ram_mem1_76_13, p_wishbone_bd_ram_mem1_76_14,
         p_wishbone_bd_ram_mem1_76_15, p_wishbone_bd_ram_mem1_77_8,
         p_wishbone_bd_ram_mem1_77_9, p_wishbone_bd_ram_mem1_77_10,
         p_wishbone_bd_ram_mem1_77_11, p_wishbone_bd_ram_mem1_77_12,
         p_wishbone_bd_ram_mem1_77_13, p_wishbone_bd_ram_mem1_77_14,
         p_wishbone_bd_ram_mem1_77_15, p_wishbone_bd_ram_mem1_78_8,
         p_wishbone_bd_ram_mem1_78_9, p_wishbone_bd_ram_mem1_78_10,
         p_wishbone_bd_ram_mem1_78_11, p_wishbone_bd_ram_mem1_78_12,
         p_wishbone_bd_ram_mem1_78_13, p_wishbone_bd_ram_mem1_78_14,
         p_wishbone_bd_ram_mem1_78_15, p_wishbone_bd_ram_mem1_79_8,
         p_wishbone_bd_ram_mem1_79_9, p_wishbone_bd_ram_mem1_79_10,
         p_wishbone_bd_ram_mem1_79_11, p_wishbone_bd_ram_mem1_79_12,
         p_wishbone_bd_ram_mem1_79_13, p_wishbone_bd_ram_mem1_79_14,
         p_wishbone_bd_ram_mem1_79_15, p_wishbone_bd_ram_mem1_80_8,
         p_wishbone_bd_ram_mem1_80_9, p_wishbone_bd_ram_mem1_80_10,
         p_wishbone_bd_ram_mem1_80_11, p_wishbone_bd_ram_mem1_80_12,
         p_wishbone_bd_ram_mem1_80_13, p_wishbone_bd_ram_mem1_80_14,
         p_wishbone_bd_ram_mem1_80_15, p_wishbone_bd_ram_mem1_81_8,
         p_wishbone_bd_ram_mem1_81_9, p_wishbone_bd_ram_mem1_81_10,
         p_wishbone_bd_ram_mem1_81_11, p_wishbone_bd_ram_mem1_81_12,
         p_wishbone_bd_ram_mem1_81_13, p_wishbone_bd_ram_mem1_81_14,
         p_wishbone_bd_ram_mem1_81_15, p_wishbone_bd_ram_mem1_82_8,
         p_wishbone_bd_ram_mem1_82_9, p_wishbone_bd_ram_mem1_82_10,
         p_wishbone_bd_ram_mem1_82_11, p_wishbone_bd_ram_mem1_82_12,
         p_wishbone_bd_ram_mem1_82_13, p_wishbone_bd_ram_mem1_82_14,
         p_wishbone_bd_ram_mem1_82_15, p_wishbone_bd_ram_mem1_83_8,
         p_wishbone_bd_ram_mem1_83_9, p_wishbone_bd_ram_mem1_83_10,
         p_wishbone_bd_ram_mem1_83_11, p_wishbone_bd_ram_mem1_83_12,
         p_wishbone_bd_ram_mem1_83_13, p_wishbone_bd_ram_mem1_83_14,
         p_wishbone_bd_ram_mem1_83_15, p_wishbone_bd_ram_mem1_84_8,
         p_wishbone_bd_ram_mem1_84_9, p_wishbone_bd_ram_mem1_84_10,
         p_wishbone_bd_ram_mem1_84_11, p_wishbone_bd_ram_mem1_84_12,
         p_wishbone_bd_ram_mem1_84_13, p_wishbone_bd_ram_mem1_84_14,
         p_wishbone_bd_ram_mem1_84_15, p_wishbone_bd_ram_mem1_85_8,
         p_wishbone_bd_ram_mem1_85_9, p_wishbone_bd_ram_mem1_85_10,
         p_wishbone_bd_ram_mem1_85_11, p_wishbone_bd_ram_mem1_85_12,
         p_wishbone_bd_ram_mem1_85_13, p_wishbone_bd_ram_mem1_85_14,
         p_wishbone_bd_ram_mem1_85_15, p_wishbone_bd_ram_mem1_86_8,
         p_wishbone_bd_ram_mem1_86_9, p_wishbone_bd_ram_mem1_86_10,
         p_wishbone_bd_ram_mem1_86_11, p_wishbone_bd_ram_mem1_86_12,
         p_wishbone_bd_ram_mem1_86_13, p_wishbone_bd_ram_mem1_86_14,
         p_wishbone_bd_ram_mem1_86_15, p_wishbone_bd_ram_mem1_87_8,
         p_wishbone_bd_ram_mem1_87_9, p_wishbone_bd_ram_mem1_87_10,
         p_wishbone_bd_ram_mem1_87_11, p_wishbone_bd_ram_mem1_87_12,
         p_wishbone_bd_ram_mem1_87_13, p_wishbone_bd_ram_mem1_87_14,
         p_wishbone_bd_ram_mem1_87_15, p_wishbone_bd_ram_mem1_88_8,
         p_wishbone_bd_ram_mem1_88_9, p_wishbone_bd_ram_mem1_88_10,
         p_wishbone_bd_ram_mem1_88_11, p_wishbone_bd_ram_mem1_88_12,
         p_wishbone_bd_ram_mem1_88_13, p_wishbone_bd_ram_mem1_88_14,
         p_wishbone_bd_ram_mem1_88_15, p_wishbone_bd_ram_mem1_89_8,
         p_wishbone_bd_ram_mem1_89_9, p_wishbone_bd_ram_mem1_89_10,
         p_wishbone_bd_ram_mem1_89_11, p_wishbone_bd_ram_mem1_89_12,
         p_wishbone_bd_ram_mem1_89_13, p_wishbone_bd_ram_mem1_89_14,
         p_wishbone_bd_ram_mem1_89_15, p_wishbone_bd_ram_mem1_90_8,
         p_wishbone_bd_ram_mem1_90_9, p_wishbone_bd_ram_mem1_90_10,
         p_wishbone_bd_ram_mem1_90_11, p_wishbone_bd_ram_mem1_90_12,
         p_wishbone_bd_ram_mem1_90_13, p_wishbone_bd_ram_mem1_90_14,
         p_wishbone_bd_ram_mem1_90_15, p_wishbone_bd_ram_mem1_91_8,
         p_wishbone_bd_ram_mem1_91_9, p_wishbone_bd_ram_mem1_91_10,
         p_wishbone_bd_ram_mem1_91_11, p_wishbone_bd_ram_mem1_91_12,
         p_wishbone_bd_ram_mem1_91_13, p_wishbone_bd_ram_mem1_91_14,
         p_wishbone_bd_ram_mem1_91_15, p_wishbone_bd_ram_mem1_92_8,
         p_wishbone_bd_ram_mem1_92_9, p_wishbone_bd_ram_mem1_92_10,
         p_wishbone_bd_ram_mem1_92_11, p_wishbone_bd_ram_mem1_92_12,
         p_wishbone_bd_ram_mem1_92_13, p_wishbone_bd_ram_mem1_92_14,
         p_wishbone_bd_ram_mem1_92_15, p_wishbone_bd_ram_mem1_93_8,
         p_wishbone_bd_ram_mem1_93_9, p_wishbone_bd_ram_mem1_93_10,
         p_wishbone_bd_ram_mem1_93_11, p_wishbone_bd_ram_mem1_93_12,
         p_wishbone_bd_ram_mem1_93_13, p_wishbone_bd_ram_mem1_93_14,
         p_wishbone_bd_ram_mem1_93_15, p_wishbone_bd_ram_mem1_94_8,
         p_wishbone_bd_ram_mem1_94_9, p_wishbone_bd_ram_mem1_94_10,
         p_wishbone_bd_ram_mem1_94_11, p_wishbone_bd_ram_mem1_94_12,
         p_wishbone_bd_ram_mem1_94_13, p_wishbone_bd_ram_mem1_94_14,
         p_wishbone_bd_ram_mem1_94_15, p_wishbone_bd_ram_mem1_95_8,
         p_wishbone_bd_ram_mem1_95_9, p_wishbone_bd_ram_mem1_95_10,
         p_wishbone_bd_ram_mem1_95_11, p_wishbone_bd_ram_mem1_95_12,
         p_wishbone_bd_ram_mem1_95_13, p_wishbone_bd_ram_mem1_95_14,
         p_wishbone_bd_ram_mem1_95_15, p_wishbone_bd_ram_mem1_96_8,
         p_wishbone_bd_ram_mem1_96_9, p_wishbone_bd_ram_mem1_96_10,
         p_wishbone_bd_ram_mem1_96_11, p_wishbone_bd_ram_mem1_96_12,
         p_wishbone_bd_ram_mem1_96_13, p_wishbone_bd_ram_mem1_96_14,
         p_wishbone_bd_ram_mem1_96_15, p_wishbone_bd_ram_mem1_97_8,
         p_wishbone_bd_ram_mem1_97_9, p_wishbone_bd_ram_mem1_97_10,
         p_wishbone_bd_ram_mem1_97_11, p_wishbone_bd_ram_mem1_97_12,
         p_wishbone_bd_ram_mem1_97_13, p_wishbone_bd_ram_mem1_97_14,
         p_wishbone_bd_ram_mem1_97_15, p_wishbone_bd_ram_mem1_98_8,
         p_wishbone_bd_ram_mem1_98_9, p_wishbone_bd_ram_mem1_98_10,
         p_wishbone_bd_ram_mem1_98_11, p_wishbone_bd_ram_mem1_98_12,
         p_wishbone_bd_ram_mem1_98_13, p_wishbone_bd_ram_mem1_98_14,
         p_wishbone_bd_ram_mem1_98_15, p_wishbone_bd_ram_mem1_99_8,
         p_wishbone_bd_ram_mem1_99_9, p_wishbone_bd_ram_mem1_99_10,
         p_wishbone_bd_ram_mem1_99_11, p_wishbone_bd_ram_mem1_99_12,
         p_wishbone_bd_ram_mem1_99_13, p_wishbone_bd_ram_mem1_99_14,
         p_wishbone_bd_ram_mem1_99_15, p_wishbone_bd_ram_mem1_100_8,
         p_wishbone_bd_ram_mem1_100_9, p_wishbone_bd_ram_mem1_100_10,
         p_wishbone_bd_ram_mem1_100_11, p_wishbone_bd_ram_mem1_100_12,
         p_wishbone_bd_ram_mem1_100_13, p_wishbone_bd_ram_mem1_100_14,
         p_wishbone_bd_ram_mem1_100_15, p_wishbone_bd_ram_mem1_101_8,
         p_wishbone_bd_ram_mem1_101_9, p_wishbone_bd_ram_mem1_101_10,
         p_wishbone_bd_ram_mem1_101_11, p_wishbone_bd_ram_mem1_101_12,
         p_wishbone_bd_ram_mem1_101_13, p_wishbone_bd_ram_mem1_101_14,
         p_wishbone_bd_ram_mem1_101_15, p_wishbone_bd_ram_mem1_102_8,
         p_wishbone_bd_ram_mem1_102_9, p_wishbone_bd_ram_mem1_102_10,
         p_wishbone_bd_ram_mem1_102_11, p_wishbone_bd_ram_mem1_102_12,
         p_wishbone_bd_ram_mem1_102_13, p_wishbone_bd_ram_mem1_102_14,
         p_wishbone_bd_ram_mem1_102_15, p_wishbone_bd_ram_mem1_103_8,
         p_wishbone_bd_ram_mem1_103_9, p_wishbone_bd_ram_mem1_103_10,
         p_wishbone_bd_ram_mem1_103_11, p_wishbone_bd_ram_mem1_103_12,
         p_wishbone_bd_ram_mem1_103_13, p_wishbone_bd_ram_mem1_103_14,
         p_wishbone_bd_ram_mem1_103_15, p_wishbone_bd_ram_mem1_104_8,
         p_wishbone_bd_ram_mem1_104_9, p_wishbone_bd_ram_mem1_104_10,
         p_wishbone_bd_ram_mem1_104_11, p_wishbone_bd_ram_mem1_104_12,
         p_wishbone_bd_ram_mem1_104_13, p_wishbone_bd_ram_mem1_104_14,
         p_wishbone_bd_ram_mem1_104_15, p_wishbone_bd_ram_mem1_105_8,
         p_wishbone_bd_ram_mem1_105_9, p_wishbone_bd_ram_mem1_105_10,
         p_wishbone_bd_ram_mem1_105_11, p_wishbone_bd_ram_mem1_105_12,
         p_wishbone_bd_ram_mem1_105_13, p_wishbone_bd_ram_mem1_105_14,
         p_wishbone_bd_ram_mem1_105_15, p_wishbone_bd_ram_mem1_106_8,
         p_wishbone_bd_ram_mem1_106_9, p_wishbone_bd_ram_mem1_106_10,
         p_wishbone_bd_ram_mem1_106_11, p_wishbone_bd_ram_mem1_106_12,
         p_wishbone_bd_ram_mem1_106_13, p_wishbone_bd_ram_mem1_106_14,
         p_wishbone_bd_ram_mem1_106_15, p_wishbone_bd_ram_mem1_107_8,
         p_wishbone_bd_ram_mem1_107_9, p_wishbone_bd_ram_mem1_107_10,
         p_wishbone_bd_ram_mem1_107_11, p_wishbone_bd_ram_mem1_107_12,
         p_wishbone_bd_ram_mem1_107_13, p_wishbone_bd_ram_mem1_107_14,
         p_wishbone_bd_ram_mem1_107_15, p_wishbone_bd_ram_mem1_108_8,
         p_wishbone_bd_ram_mem1_108_9, p_wishbone_bd_ram_mem1_108_10,
         p_wishbone_bd_ram_mem1_108_11, p_wishbone_bd_ram_mem1_108_12,
         p_wishbone_bd_ram_mem1_108_13, p_wishbone_bd_ram_mem1_108_14,
         p_wishbone_bd_ram_mem1_108_15, p_wishbone_bd_ram_mem1_109_8,
         p_wishbone_bd_ram_mem1_109_9, p_wishbone_bd_ram_mem1_109_10,
         p_wishbone_bd_ram_mem1_109_11, p_wishbone_bd_ram_mem1_109_12,
         p_wishbone_bd_ram_mem1_109_13, p_wishbone_bd_ram_mem1_109_14,
         p_wishbone_bd_ram_mem1_109_15, p_wishbone_bd_ram_mem1_110_8,
         p_wishbone_bd_ram_mem1_110_9, p_wishbone_bd_ram_mem1_110_10,
         p_wishbone_bd_ram_mem1_110_11, p_wishbone_bd_ram_mem1_110_12,
         p_wishbone_bd_ram_mem1_110_13, p_wishbone_bd_ram_mem1_110_14,
         p_wishbone_bd_ram_mem1_110_15, p_wishbone_bd_ram_mem1_111_8,
         p_wishbone_bd_ram_mem1_111_9, p_wishbone_bd_ram_mem1_111_10,
         p_wishbone_bd_ram_mem1_111_11, p_wishbone_bd_ram_mem1_111_12,
         p_wishbone_bd_ram_mem1_111_13, p_wishbone_bd_ram_mem1_111_14,
         p_wishbone_bd_ram_mem1_111_15, p_wishbone_bd_ram_mem1_112_8,
         p_wishbone_bd_ram_mem1_112_9, p_wishbone_bd_ram_mem1_112_10,
         p_wishbone_bd_ram_mem1_112_11, p_wishbone_bd_ram_mem1_112_12,
         p_wishbone_bd_ram_mem1_112_13, p_wishbone_bd_ram_mem1_112_14,
         p_wishbone_bd_ram_mem1_112_15, p_wishbone_bd_ram_mem1_113_8,
         p_wishbone_bd_ram_mem1_113_9, p_wishbone_bd_ram_mem1_113_10,
         p_wishbone_bd_ram_mem1_113_11, p_wishbone_bd_ram_mem1_113_12,
         p_wishbone_bd_ram_mem1_113_13, p_wishbone_bd_ram_mem1_113_14,
         p_wishbone_bd_ram_mem1_113_15, p_wishbone_bd_ram_mem1_114_8,
         p_wishbone_bd_ram_mem1_114_9, p_wishbone_bd_ram_mem1_114_10,
         p_wishbone_bd_ram_mem1_114_11, p_wishbone_bd_ram_mem1_114_12,
         p_wishbone_bd_ram_mem1_114_13, p_wishbone_bd_ram_mem1_114_14,
         p_wishbone_bd_ram_mem1_114_15, p_wishbone_bd_ram_mem1_115_8,
         p_wishbone_bd_ram_mem1_115_9, p_wishbone_bd_ram_mem1_115_10,
         p_wishbone_bd_ram_mem1_115_11, p_wishbone_bd_ram_mem1_115_12,
         p_wishbone_bd_ram_mem1_115_13, p_wishbone_bd_ram_mem1_115_14,
         p_wishbone_bd_ram_mem1_115_15, p_wishbone_bd_ram_mem1_116_8,
         p_wishbone_bd_ram_mem1_116_9, p_wishbone_bd_ram_mem1_116_10,
         p_wishbone_bd_ram_mem1_116_11, p_wishbone_bd_ram_mem1_116_12,
         p_wishbone_bd_ram_mem1_116_13, p_wishbone_bd_ram_mem1_116_14,
         p_wishbone_bd_ram_mem1_116_15, p_wishbone_bd_ram_mem1_117_8,
         p_wishbone_bd_ram_mem1_117_9, p_wishbone_bd_ram_mem1_117_10,
         p_wishbone_bd_ram_mem1_117_11, p_wishbone_bd_ram_mem1_117_12,
         p_wishbone_bd_ram_mem1_117_13, p_wishbone_bd_ram_mem1_117_14,
         p_wishbone_bd_ram_mem1_117_15, p_wishbone_bd_ram_mem1_118_8,
         p_wishbone_bd_ram_mem1_118_9, p_wishbone_bd_ram_mem1_118_10,
         p_wishbone_bd_ram_mem1_118_11, p_wishbone_bd_ram_mem1_118_12,
         p_wishbone_bd_ram_mem1_118_13, p_wishbone_bd_ram_mem1_118_14,
         p_wishbone_bd_ram_mem1_118_15, p_wishbone_bd_ram_mem1_119_8,
         p_wishbone_bd_ram_mem1_119_9, p_wishbone_bd_ram_mem1_119_10,
         p_wishbone_bd_ram_mem1_119_11, p_wishbone_bd_ram_mem1_119_12,
         p_wishbone_bd_ram_mem1_119_13, p_wishbone_bd_ram_mem1_119_14,
         p_wishbone_bd_ram_mem1_119_15, p_wishbone_bd_ram_mem1_120_8,
         p_wishbone_bd_ram_mem1_120_9, p_wishbone_bd_ram_mem1_120_10,
         p_wishbone_bd_ram_mem1_120_11, p_wishbone_bd_ram_mem1_120_12,
         p_wishbone_bd_ram_mem1_120_13, p_wishbone_bd_ram_mem1_120_14,
         p_wishbone_bd_ram_mem1_120_15, p_wishbone_bd_ram_mem1_121_8,
         p_wishbone_bd_ram_mem1_121_9, p_wishbone_bd_ram_mem1_121_10,
         p_wishbone_bd_ram_mem1_121_11, p_wishbone_bd_ram_mem1_121_12,
         p_wishbone_bd_ram_mem1_121_13, p_wishbone_bd_ram_mem1_121_14,
         p_wishbone_bd_ram_mem1_121_15, p_wishbone_bd_ram_mem1_122_8,
         p_wishbone_bd_ram_mem1_122_9, p_wishbone_bd_ram_mem1_122_10,
         p_wishbone_bd_ram_mem1_122_11, p_wishbone_bd_ram_mem1_122_12,
         p_wishbone_bd_ram_mem1_122_13, p_wishbone_bd_ram_mem1_122_14,
         p_wishbone_bd_ram_mem1_122_15, p_wishbone_bd_ram_mem1_123_8,
         p_wishbone_bd_ram_mem1_123_9, p_wishbone_bd_ram_mem1_123_10,
         p_wishbone_bd_ram_mem1_123_11, p_wishbone_bd_ram_mem1_123_12,
         p_wishbone_bd_ram_mem1_123_13, p_wishbone_bd_ram_mem1_123_14,
         p_wishbone_bd_ram_mem1_123_15, p_wishbone_bd_ram_mem1_124_8,
         p_wishbone_bd_ram_mem1_124_9, p_wishbone_bd_ram_mem1_124_10,
         p_wishbone_bd_ram_mem1_124_11, p_wishbone_bd_ram_mem1_124_12,
         p_wishbone_bd_ram_mem1_124_13, p_wishbone_bd_ram_mem1_124_14,
         p_wishbone_bd_ram_mem1_124_15, p_wishbone_bd_ram_mem1_125_8,
         p_wishbone_bd_ram_mem1_125_9, p_wishbone_bd_ram_mem1_125_10,
         p_wishbone_bd_ram_mem1_125_11, p_wishbone_bd_ram_mem1_125_12,
         p_wishbone_bd_ram_mem1_125_13, p_wishbone_bd_ram_mem1_125_14,
         p_wishbone_bd_ram_mem1_125_15, p_wishbone_bd_ram_mem1_126_8,
         p_wishbone_bd_ram_mem1_126_9, p_wishbone_bd_ram_mem1_126_10,
         p_wishbone_bd_ram_mem1_126_11, p_wishbone_bd_ram_mem1_126_12,
         p_wishbone_bd_ram_mem1_126_13, p_wishbone_bd_ram_mem1_126_14,
         p_wishbone_bd_ram_mem1_126_15, p_wishbone_bd_ram_mem1_127_8,
         p_wishbone_bd_ram_mem1_127_9, p_wishbone_bd_ram_mem1_127_10,
         p_wishbone_bd_ram_mem1_127_11, p_wishbone_bd_ram_mem1_127_12,
         p_wishbone_bd_ram_mem1_127_13, p_wishbone_bd_ram_mem1_127_14,
         p_wishbone_bd_ram_mem1_127_15, p_wishbone_bd_ram_mem1_128_8,
         p_wishbone_bd_ram_mem1_128_9, p_wishbone_bd_ram_mem1_128_10,
         p_wishbone_bd_ram_mem1_128_11, p_wishbone_bd_ram_mem1_128_12,
         p_wishbone_bd_ram_mem1_128_13, p_wishbone_bd_ram_mem1_128_14,
         p_wishbone_bd_ram_mem1_128_15, p_wishbone_bd_ram_mem1_129_8,
         p_wishbone_bd_ram_mem1_129_9, p_wishbone_bd_ram_mem1_129_10,
         p_wishbone_bd_ram_mem1_129_11, p_wishbone_bd_ram_mem1_129_12,
         p_wishbone_bd_ram_mem1_129_13, p_wishbone_bd_ram_mem1_129_14,
         p_wishbone_bd_ram_mem1_129_15, p_wishbone_bd_ram_mem1_130_8,
         p_wishbone_bd_ram_mem1_130_9, p_wishbone_bd_ram_mem1_130_10,
         p_wishbone_bd_ram_mem1_130_11, p_wishbone_bd_ram_mem1_130_12,
         p_wishbone_bd_ram_mem1_130_13, p_wishbone_bd_ram_mem1_130_14,
         p_wishbone_bd_ram_mem1_130_15, p_wishbone_bd_ram_mem1_131_8,
         p_wishbone_bd_ram_mem1_131_9, p_wishbone_bd_ram_mem1_131_10,
         p_wishbone_bd_ram_mem1_131_11, p_wishbone_bd_ram_mem1_131_12,
         p_wishbone_bd_ram_mem1_131_13, p_wishbone_bd_ram_mem1_131_14,
         p_wishbone_bd_ram_mem1_131_15, p_wishbone_bd_ram_mem1_132_8,
         p_wishbone_bd_ram_mem1_132_9, p_wishbone_bd_ram_mem1_132_10,
         p_wishbone_bd_ram_mem1_132_11, p_wishbone_bd_ram_mem1_132_12,
         p_wishbone_bd_ram_mem1_132_13, p_wishbone_bd_ram_mem1_132_14,
         p_wishbone_bd_ram_mem1_132_15, p_wishbone_bd_ram_mem1_133_8,
         p_wishbone_bd_ram_mem1_133_9, p_wishbone_bd_ram_mem1_133_10,
         p_wishbone_bd_ram_mem1_133_11, p_wishbone_bd_ram_mem1_133_12,
         p_wishbone_bd_ram_mem1_133_13, p_wishbone_bd_ram_mem1_133_14,
         p_wishbone_bd_ram_mem1_133_15, p_wishbone_bd_ram_mem1_134_8,
         p_wishbone_bd_ram_mem1_134_9, p_wishbone_bd_ram_mem1_134_10,
         p_wishbone_bd_ram_mem1_134_11, p_wishbone_bd_ram_mem1_134_12,
         p_wishbone_bd_ram_mem1_134_13, p_wishbone_bd_ram_mem1_134_14,
         p_wishbone_bd_ram_mem1_134_15, p_wishbone_bd_ram_mem1_135_8,
         p_wishbone_bd_ram_mem1_135_9, p_wishbone_bd_ram_mem1_135_10,
         p_wishbone_bd_ram_mem1_135_11, p_wishbone_bd_ram_mem1_135_12,
         p_wishbone_bd_ram_mem1_135_13, p_wishbone_bd_ram_mem1_135_14,
         p_wishbone_bd_ram_mem1_135_15, p_wishbone_bd_ram_mem1_136_8,
         p_wishbone_bd_ram_mem1_136_9, p_wishbone_bd_ram_mem1_136_10,
         p_wishbone_bd_ram_mem1_136_11, p_wishbone_bd_ram_mem1_136_12,
         p_wishbone_bd_ram_mem1_136_13, p_wishbone_bd_ram_mem1_136_14,
         p_wishbone_bd_ram_mem1_136_15, p_wishbone_bd_ram_mem1_137_8,
         p_wishbone_bd_ram_mem1_137_9, p_wishbone_bd_ram_mem1_137_10,
         p_wishbone_bd_ram_mem1_137_11, p_wishbone_bd_ram_mem1_137_12,
         p_wishbone_bd_ram_mem1_137_13, p_wishbone_bd_ram_mem1_137_14,
         p_wishbone_bd_ram_mem1_137_15, p_wishbone_bd_ram_mem1_138_8,
         p_wishbone_bd_ram_mem1_138_9, p_wishbone_bd_ram_mem1_138_10,
         p_wishbone_bd_ram_mem1_138_11, p_wishbone_bd_ram_mem1_138_12,
         p_wishbone_bd_ram_mem1_138_13, p_wishbone_bd_ram_mem1_138_14,
         p_wishbone_bd_ram_mem1_138_15, p_wishbone_bd_ram_mem1_139_8,
         p_wishbone_bd_ram_mem1_139_9, p_wishbone_bd_ram_mem1_139_10,
         p_wishbone_bd_ram_mem1_139_11, p_wishbone_bd_ram_mem1_139_12,
         p_wishbone_bd_ram_mem1_139_13, p_wishbone_bd_ram_mem1_139_14,
         p_wishbone_bd_ram_mem1_139_15, p_wishbone_bd_ram_mem1_140_8,
         p_wishbone_bd_ram_mem1_140_9, p_wishbone_bd_ram_mem1_140_10,
         p_wishbone_bd_ram_mem1_140_11, p_wishbone_bd_ram_mem1_140_12,
         p_wishbone_bd_ram_mem1_140_13, p_wishbone_bd_ram_mem1_140_14,
         p_wishbone_bd_ram_mem1_140_15, p_wishbone_bd_ram_mem1_141_8,
         p_wishbone_bd_ram_mem1_141_9, p_wishbone_bd_ram_mem1_141_10,
         p_wishbone_bd_ram_mem1_141_11, p_wishbone_bd_ram_mem1_141_12,
         p_wishbone_bd_ram_mem1_141_13, p_wishbone_bd_ram_mem1_141_14,
         p_wishbone_bd_ram_mem1_141_15, p_wishbone_bd_ram_mem1_142_8,
         p_wishbone_bd_ram_mem1_142_9, p_wishbone_bd_ram_mem1_142_10,
         p_wishbone_bd_ram_mem1_142_11, p_wishbone_bd_ram_mem1_142_12,
         p_wishbone_bd_ram_mem1_142_13, p_wishbone_bd_ram_mem1_142_14,
         p_wishbone_bd_ram_mem1_142_15, p_wishbone_bd_ram_mem1_143_8,
         p_wishbone_bd_ram_mem1_143_9, p_wishbone_bd_ram_mem1_143_10,
         p_wishbone_bd_ram_mem1_143_11, p_wishbone_bd_ram_mem1_143_12,
         p_wishbone_bd_ram_mem1_143_13, p_wishbone_bd_ram_mem1_143_14,
         p_wishbone_bd_ram_mem1_143_15, p_wishbone_bd_ram_mem1_144_8,
         p_wishbone_bd_ram_mem1_144_9, p_wishbone_bd_ram_mem1_144_10,
         p_wishbone_bd_ram_mem1_144_11, p_wishbone_bd_ram_mem1_144_12,
         p_wishbone_bd_ram_mem1_144_13, p_wishbone_bd_ram_mem1_144_14,
         p_wishbone_bd_ram_mem1_144_15, p_wishbone_bd_ram_mem1_145_8,
         p_wishbone_bd_ram_mem1_145_9, p_wishbone_bd_ram_mem1_145_10,
         p_wishbone_bd_ram_mem1_145_11, p_wishbone_bd_ram_mem1_145_12,
         p_wishbone_bd_ram_mem1_145_13, p_wishbone_bd_ram_mem1_145_14,
         p_wishbone_bd_ram_mem1_145_15, p_wishbone_bd_ram_mem1_146_8,
         p_wishbone_bd_ram_mem1_146_9, p_wishbone_bd_ram_mem1_146_10,
         p_wishbone_bd_ram_mem1_146_11, p_wishbone_bd_ram_mem1_146_12,
         p_wishbone_bd_ram_mem1_146_13, p_wishbone_bd_ram_mem1_146_14,
         p_wishbone_bd_ram_mem1_146_15, p_wishbone_bd_ram_mem1_147_8,
         p_wishbone_bd_ram_mem1_147_9, p_wishbone_bd_ram_mem1_147_10,
         p_wishbone_bd_ram_mem1_147_11, p_wishbone_bd_ram_mem1_147_12,
         p_wishbone_bd_ram_mem1_147_13, p_wishbone_bd_ram_mem1_147_14,
         p_wishbone_bd_ram_mem1_147_15, p_wishbone_bd_ram_mem1_148_8,
         p_wishbone_bd_ram_mem1_148_9, p_wishbone_bd_ram_mem1_148_10,
         p_wishbone_bd_ram_mem1_148_11, p_wishbone_bd_ram_mem1_148_12,
         p_wishbone_bd_ram_mem1_148_13, p_wishbone_bd_ram_mem1_148_14,
         p_wishbone_bd_ram_mem1_148_15, p_wishbone_bd_ram_mem1_149_8,
         p_wishbone_bd_ram_mem1_149_9, p_wishbone_bd_ram_mem1_149_10,
         p_wishbone_bd_ram_mem1_149_11, p_wishbone_bd_ram_mem1_149_12,
         p_wishbone_bd_ram_mem1_149_13, p_wishbone_bd_ram_mem1_149_14,
         p_wishbone_bd_ram_mem1_149_15, p_wishbone_bd_ram_mem1_150_8,
         p_wishbone_bd_ram_mem1_150_9, p_wishbone_bd_ram_mem1_150_10,
         p_wishbone_bd_ram_mem1_150_11, p_wishbone_bd_ram_mem1_150_12,
         p_wishbone_bd_ram_mem1_150_13, p_wishbone_bd_ram_mem1_150_14,
         p_wishbone_bd_ram_mem1_150_15, p_wishbone_bd_ram_mem1_151_8,
         p_wishbone_bd_ram_mem1_151_9, p_wishbone_bd_ram_mem1_151_10,
         p_wishbone_bd_ram_mem1_151_11, p_wishbone_bd_ram_mem1_151_12,
         p_wishbone_bd_ram_mem1_151_13, p_wishbone_bd_ram_mem1_151_14,
         p_wishbone_bd_ram_mem1_151_15, p_wishbone_bd_ram_mem1_152_8,
         p_wishbone_bd_ram_mem1_152_9, p_wishbone_bd_ram_mem1_152_10,
         p_wishbone_bd_ram_mem1_152_11, p_wishbone_bd_ram_mem1_152_12,
         p_wishbone_bd_ram_mem1_152_13, p_wishbone_bd_ram_mem1_152_14,
         p_wishbone_bd_ram_mem1_152_15, p_wishbone_bd_ram_mem1_153_8,
         p_wishbone_bd_ram_mem1_153_9, p_wishbone_bd_ram_mem1_153_10,
         p_wishbone_bd_ram_mem1_153_11, p_wishbone_bd_ram_mem1_153_12,
         p_wishbone_bd_ram_mem1_153_13, p_wishbone_bd_ram_mem1_153_14,
         p_wishbone_bd_ram_mem1_153_15, p_wishbone_bd_ram_mem1_154_8,
         p_wishbone_bd_ram_mem1_154_9, p_wishbone_bd_ram_mem1_154_10,
         p_wishbone_bd_ram_mem1_154_11, p_wishbone_bd_ram_mem1_154_12,
         p_wishbone_bd_ram_mem1_154_13, p_wishbone_bd_ram_mem1_154_14,
         p_wishbone_bd_ram_mem1_154_15, p_wishbone_bd_ram_mem1_155_8,
         p_wishbone_bd_ram_mem1_155_9, p_wishbone_bd_ram_mem1_155_10,
         p_wishbone_bd_ram_mem1_155_11, p_wishbone_bd_ram_mem1_155_12,
         p_wishbone_bd_ram_mem1_155_13, p_wishbone_bd_ram_mem1_155_14,
         p_wishbone_bd_ram_mem1_155_15, p_wishbone_bd_ram_mem1_156_8,
         p_wishbone_bd_ram_mem1_156_9, p_wishbone_bd_ram_mem1_156_10,
         p_wishbone_bd_ram_mem1_156_11, p_wishbone_bd_ram_mem1_156_12,
         p_wishbone_bd_ram_mem1_156_13, p_wishbone_bd_ram_mem1_156_14,
         p_wishbone_bd_ram_mem1_156_15, p_wishbone_bd_ram_mem1_157_8,
         p_wishbone_bd_ram_mem1_157_9, p_wishbone_bd_ram_mem1_157_10,
         p_wishbone_bd_ram_mem1_157_11, p_wishbone_bd_ram_mem1_157_12,
         p_wishbone_bd_ram_mem1_157_13, p_wishbone_bd_ram_mem1_157_14,
         p_wishbone_bd_ram_mem1_157_15, p_wishbone_bd_ram_mem1_158_8,
         p_wishbone_bd_ram_mem1_158_9, p_wishbone_bd_ram_mem1_158_10,
         p_wishbone_bd_ram_mem1_158_11, p_wishbone_bd_ram_mem1_158_12,
         p_wishbone_bd_ram_mem1_158_13, p_wishbone_bd_ram_mem1_158_14,
         p_wishbone_bd_ram_mem1_158_15, p_wishbone_bd_ram_mem1_159_8,
         p_wishbone_bd_ram_mem1_159_9, p_wishbone_bd_ram_mem1_159_10,
         p_wishbone_bd_ram_mem1_159_11, p_wishbone_bd_ram_mem1_159_12,
         p_wishbone_bd_ram_mem1_159_13, p_wishbone_bd_ram_mem1_159_14,
         p_wishbone_bd_ram_mem1_159_15, p_wishbone_bd_ram_mem1_160_8,
         p_wishbone_bd_ram_mem1_160_9, p_wishbone_bd_ram_mem1_160_10,
         p_wishbone_bd_ram_mem1_160_11, p_wishbone_bd_ram_mem1_160_12,
         p_wishbone_bd_ram_mem1_160_13, p_wishbone_bd_ram_mem1_160_14,
         p_wishbone_bd_ram_mem1_160_15, p_wishbone_bd_ram_mem1_161_8,
         p_wishbone_bd_ram_mem1_161_9, p_wishbone_bd_ram_mem1_161_10,
         p_wishbone_bd_ram_mem1_161_11, p_wishbone_bd_ram_mem1_161_12,
         p_wishbone_bd_ram_mem1_161_13, p_wishbone_bd_ram_mem1_161_14,
         p_wishbone_bd_ram_mem1_161_15, p_wishbone_bd_ram_mem1_162_8,
         p_wishbone_bd_ram_mem1_162_9, p_wishbone_bd_ram_mem1_162_10,
         p_wishbone_bd_ram_mem1_162_11, p_wishbone_bd_ram_mem1_162_12,
         p_wishbone_bd_ram_mem1_162_13, p_wishbone_bd_ram_mem1_162_14,
         p_wishbone_bd_ram_mem1_162_15, p_wishbone_bd_ram_mem1_163_8,
         p_wishbone_bd_ram_mem1_163_9, p_wishbone_bd_ram_mem1_163_10,
         p_wishbone_bd_ram_mem1_163_11, p_wishbone_bd_ram_mem1_163_12,
         p_wishbone_bd_ram_mem1_163_13, p_wishbone_bd_ram_mem1_163_14,
         p_wishbone_bd_ram_mem1_163_15, p_wishbone_bd_ram_mem1_164_8,
         p_wishbone_bd_ram_mem1_164_9, p_wishbone_bd_ram_mem1_164_10,
         p_wishbone_bd_ram_mem1_164_11, p_wishbone_bd_ram_mem1_164_12,
         p_wishbone_bd_ram_mem1_164_13, p_wishbone_bd_ram_mem1_164_14,
         p_wishbone_bd_ram_mem1_164_15, p_wishbone_bd_ram_mem1_165_8,
         p_wishbone_bd_ram_mem1_165_9, p_wishbone_bd_ram_mem1_165_10,
         p_wishbone_bd_ram_mem1_165_11, p_wishbone_bd_ram_mem1_165_12,
         p_wishbone_bd_ram_mem1_165_13, p_wishbone_bd_ram_mem1_165_14,
         p_wishbone_bd_ram_mem1_165_15, p_wishbone_bd_ram_mem1_166_8,
         p_wishbone_bd_ram_mem1_166_9, p_wishbone_bd_ram_mem1_166_10,
         p_wishbone_bd_ram_mem1_166_11, p_wishbone_bd_ram_mem1_166_12,
         p_wishbone_bd_ram_mem1_166_13, p_wishbone_bd_ram_mem1_166_14,
         p_wishbone_bd_ram_mem1_166_15, p_wishbone_bd_ram_mem1_167_8,
         p_wishbone_bd_ram_mem1_167_9, p_wishbone_bd_ram_mem1_167_10,
         p_wishbone_bd_ram_mem1_167_11, p_wishbone_bd_ram_mem1_167_12,
         p_wishbone_bd_ram_mem1_167_13, p_wishbone_bd_ram_mem1_167_14,
         p_wishbone_bd_ram_mem1_167_15, p_wishbone_bd_ram_mem1_168_8,
         p_wishbone_bd_ram_mem1_168_9, p_wishbone_bd_ram_mem1_168_10,
         p_wishbone_bd_ram_mem1_168_11, p_wishbone_bd_ram_mem1_168_12,
         p_wishbone_bd_ram_mem1_168_13, p_wishbone_bd_ram_mem1_168_14,
         p_wishbone_bd_ram_mem1_168_15, p_wishbone_bd_ram_mem1_169_8,
         p_wishbone_bd_ram_mem1_169_9, p_wishbone_bd_ram_mem1_169_10,
         p_wishbone_bd_ram_mem1_169_11, p_wishbone_bd_ram_mem1_169_12,
         p_wishbone_bd_ram_mem1_169_13, p_wishbone_bd_ram_mem1_169_14,
         p_wishbone_bd_ram_mem1_169_15, p_wishbone_bd_ram_mem1_170_8,
         p_wishbone_bd_ram_mem1_170_9, p_wishbone_bd_ram_mem1_170_10,
         p_wishbone_bd_ram_mem1_170_11, p_wishbone_bd_ram_mem1_170_12,
         p_wishbone_bd_ram_mem1_170_13, p_wishbone_bd_ram_mem1_170_14,
         p_wishbone_bd_ram_mem1_170_15, p_wishbone_bd_ram_mem1_171_8,
         p_wishbone_bd_ram_mem1_171_9, p_wishbone_bd_ram_mem1_171_10,
         p_wishbone_bd_ram_mem1_171_11, p_wishbone_bd_ram_mem1_171_12,
         p_wishbone_bd_ram_mem1_171_13, p_wishbone_bd_ram_mem1_171_14,
         p_wishbone_bd_ram_mem1_171_15, p_wishbone_bd_ram_mem1_172_8,
         p_wishbone_bd_ram_mem1_172_9, p_wishbone_bd_ram_mem1_172_10,
         p_wishbone_bd_ram_mem1_172_11, p_wishbone_bd_ram_mem1_172_12,
         p_wishbone_bd_ram_mem1_172_13, p_wishbone_bd_ram_mem1_172_14,
         p_wishbone_bd_ram_mem1_172_15, p_wishbone_bd_ram_mem1_173_8,
         p_wishbone_bd_ram_mem1_173_9, p_wishbone_bd_ram_mem1_173_10,
         p_wishbone_bd_ram_mem1_173_11, p_wishbone_bd_ram_mem1_173_12,
         p_wishbone_bd_ram_mem1_173_13, p_wishbone_bd_ram_mem1_173_14,
         p_wishbone_bd_ram_mem1_173_15, p_wishbone_bd_ram_mem1_174_8,
         p_wishbone_bd_ram_mem1_174_9, p_wishbone_bd_ram_mem1_174_10,
         p_wishbone_bd_ram_mem1_174_11, p_wishbone_bd_ram_mem1_174_12,
         p_wishbone_bd_ram_mem1_174_13, p_wishbone_bd_ram_mem1_174_14,
         p_wishbone_bd_ram_mem1_174_15, p_wishbone_bd_ram_mem1_175_8,
         p_wishbone_bd_ram_mem1_175_9, p_wishbone_bd_ram_mem1_175_10,
         p_wishbone_bd_ram_mem1_175_11, p_wishbone_bd_ram_mem1_175_12,
         p_wishbone_bd_ram_mem1_175_13, p_wishbone_bd_ram_mem1_175_14,
         p_wishbone_bd_ram_mem1_175_15, p_wishbone_bd_ram_mem1_176_8,
         p_wishbone_bd_ram_mem1_176_9, p_wishbone_bd_ram_mem1_176_10,
         p_wishbone_bd_ram_mem1_176_11, p_wishbone_bd_ram_mem1_176_12,
         p_wishbone_bd_ram_mem1_176_13, p_wishbone_bd_ram_mem1_176_14,
         p_wishbone_bd_ram_mem1_176_15, p_wishbone_bd_ram_mem1_177_8,
         p_wishbone_bd_ram_mem1_177_9, p_wishbone_bd_ram_mem1_177_10,
         p_wishbone_bd_ram_mem1_177_11, p_wishbone_bd_ram_mem1_177_12,
         p_wishbone_bd_ram_mem1_177_13, p_wishbone_bd_ram_mem1_177_14,
         p_wishbone_bd_ram_mem1_177_15, p_wishbone_bd_ram_mem1_178_8,
         p_wishbone_bd_ram_mem1_178_9, p_wishbone_bd_ram_mem1_178_10,
         p_wishbone_bd_ram_mem1_178_11, p_wishbone_bd_ram_mem1_178_12,
         p_wishbone_bd_ram_mem1_178_13, p_wishbone_bd_ram_mem1_178_14,
         p_wishbone_bd_ram_mem1_178_15, p_wishbone_bd_ram_mem1_179_8,
         p_wishbone_bd_ram_mem1_179_9, p_wishbone_bd_ram_mem1_179_10,
         p_wishbone_bd_ram_mem1_179_11, p_wishbone_bd_ram_mem1_179_12,
         p_wishbone_bd_ram_mem1_179_13, p_wishbone_bd_ram_mem1_179_14,
         p_wishbone_bd_ram_mem1_179_15, p_wishbone_bd_ram_mem1_180_8,
         p_wishbone_bd_ram_mem1_180_9, p_wishbone_bd_ram_mem1_180_10,
         p_wishbone_bd_ram_mem1_180_11, p_wishbone_bd_ram_mem1_180_12,
         p_wishbone_bd_ram_mem1_180_13, p_wishbone_bd_ram_mem1_180_14,
         p_wishbone_bd_ram_mem1_180_15, p_wishbone_bd_ram_mem1_181_8,
         p_wishbone_bd_ram_mem1_181_9, p_wishbone_bd_ram_mem1_181_10,
         p_wishbone_bd_ram_mem1_181_11, p_wishbone_bd_ram_mem1_181_12,
         p_wishbone_bd_ram_mem1_181_13, p_wishbone_bd_ram_mem1_181_14,
         p_wishbone_bd_ram_mem1_181_15, p_wishbone_bd_ram_mem1_182_8,
         p_wishbone_bd_ram_mem1_182_9, p_wishbone_bd_ram_mem1_182_10,
         p_wishbone_bd_ram_mem1_182_11, p_wishbone_bd_ram_mem1_182_12,
         p_wishbone_bd_ram_mem1_182_13, p_wishbone_bd_ram_mem1_182_14,
         p_wishbone_bd_ram_mem1_182_15, p_wishbone_bd_ram_mem1_183_8,
         p_wishbone_bd_ram_mem1_183_9, p_wishbone_bd_ram_mem1_183_10,
         p_wishbone_bd_ram_mem1_183_11, p_wishbone_bd_ram_mem1_183_12,
         p_wishbone_bd_ram_mem1_183_13, p_wishbone_bd_ram_mem1_183_14,
         p_wishbone_bd_ram_mem1_183_15, p_wishbone_bd_ram_mem1_184_8,
         p_wishbone_bd_ram_mem1_184_9, p_wishbone_bd_ram_mem1_184_10,
         p_wishbone_bd_ram_mem1_184_11, p_wishbone_bd_ram_mem1_184_12,
         p_wishbone_bd_ram_mem1_184_13, p_wishbone_bd_ram_mem1_184_14,
         p_wishbone_bd_ram_mem1_184_15, p_wishbone_bd_ram_mem1_185_8,
         p_wishbone_bd_ram_mem1_185_9, p_wishbone_bd_ram_mem1_185_10,
         p_wishbone_bd_ram_mem1_185_11, p_wishbone_bd_ram_mem1_185_12,
         p_wishbone_bd_ram_mem1_185_13, p_wishbone_bd_ram_mem1_185_14,
         p_wishbone_bd_ram_mem1_185_15, p_wishbone_bd_ram_mem1_186_8,
         p_wishbone_bd_ram_mem1_186_9, p_wishbone_bd_ram_mem1_186_10,
         p_wishbone_bd_ram_mem1_186_11, p_wishbone_bd_ram_mem1_186_12,
         p_wishbone_bd_ram_mem1_186_13, p_wishbone_bd_ram_mem1_186_14,
         p_wishbone_bd_ram_mem1_186_15, p_wishbone_bd_ram_mem1_187_8,
         p_wishbone_bd_ram_mem1_187_9, p_wishbone_bd_ram_mem1_187_10,
         p_wishbone_bd_ram_mem1_187_11, p_wishbone_bd_ram_mem1_187_12,
         p_wishbone_bd_ram_mem1_187_13, p_wishbone_bd_ram_mem1_187_14,
         p_wishbone_bd_ram_mem1_187_15, p_wishbone_bd_ram_mem1_188_8,
         p_wishbone_bd_ram_mem1_188_9, p_wishbone_bd_ram_mem1_188_10,
         p_wishbone_bd_ram_mem1_188_11, p_wishbone_bd_ram_mem1_188_12,
         p_wishbone_bd_ram_mem1_188_13, p_wishbone_bd_ram_mem1_188_14,
         p_wishbone_bd_ram_mem1_188_15, p_wishbone_bd_ram_mem1_189_8,
         p_wishbone_bd_ram_mem1_189_9, p_wishbone_bd_ram_mem1_189_10,
         p_wishbone_bd_ram_mem1_189_11, p_wishbone_bd_ram_mem1_189_12,
         p_wishbone_bd_ram_mem1_189_13, p_wishbone_bd_ram_mem1_189_14,
         p_wishbone_bd_ram_mem1_189_15, p_wishbone_bd_ram_mem1_190_8,
         p_wishbone_bd_ram_mem1_190_9, p_wishbone_bd_ram_mem1_190_10,
         p_wishbone_bd_ram_mem1_190_11, p_wishbone_bd_ram_mem1_190_12,
         p_wishbone_bd_ram_mem1_190_13, p_wishbone_bd_ram_mem1_190_14,
         p_wishbone_bd_ram_mem1_190_15, p_wishbone_bd_ram_mem1_191_8,
         p_wishbone_bd_ram_mem1_191_9, p_wishbone_bd_ram_mem1_191_10,
         p_wishbone_bd_ram_mem1_191_11, p_wishbone_bd_ram_mem1_191_12,
         p_wishbone_bd_ram_mem1_191_13, p_wishbone_bd_ram_mem1_191_14,
         p_wishbone_bd_ram_mem1_191_15, p_wishbone_bd_ram_mem1_192_8,
         p_wishbone_bd_ram_mem1_192_9, p_wishbone_bd_ram_mem1_192_10,
         p_wishbone_bd_ram_mem1_192_11, p_wishbone_bd_ram_mem1_192_12,
         p_wishbone_bd_ram_mem1_192_13, p_wishbone_bd_ram_mem1_192_14,
         p_wishbone_bd_ram_mem1_192_15, p_wishbone_bd_ram_mem1_193_8,
         p_wishbone_bd_ram_mem1_193_9, p_wishbone_bd_ram_mem1_193_10,
         p_wishbone_bd_ram_mem1_193_11, p_wishbone_bd_ram_mem1_193_12,
         p_wishbone_bd_ram_mem1_193_13, p_wishbone_bd_ram_mem1_193_14,
         p_wishbone_bd_ram_mem1_193_15, p_wishbone_bd_ram_mem1_194_8,
         p_wishbone_bd_ram_mem1_194_9, p_wishbone_bd_ram_mem1_194_10,
         p_wishbone_bd_ram_mem1_194_11, p_wishbone_bd_ram_mem1_194_12,
         p_wishbone_bd_ram_mem1_194_13, p_wishbone_bd_ram_mem1_194_14,
         p_wishbone_bd_ram_mem1_194_15, p_wishbone_bd_ram_mem1_195_8,
         p_wishbone_bd_ram_mem1_195_9, p_wishbone_bd_ram_mem1_195_10,
         p_wishbone_bd_ram_mem1_195_11, p_wishbone_bd_ram_mem1_195_12,
         p_wishbone_bd_ram_mem1_195_13, p_wishbone_bd_ram_mem1_195_14,
         p_wishbone_bd_ram_mem1_195_15, p_wishbone_bd_ram_mem1_196_8,
         p_wishbone_bd_ram_mem1_196_9, p_wishbone_bd_ram_mem1_196_10,
         p_wishbone_bd_ram_mem1_196_11, p_wishbone_bd_ram_mem1_196_12,
         p_wishbone_bd_ram_mem1_196_13, p_wishbone_bd_ram_mem1_196_14,
         p_wishbone_bd_ram_mem1_196_15, p_wishbone_bd_ram_mem1_197_8,
         p_wishbone_bd_ram_mem1_197_9, p_wishbone_bd_ram_mem1_197_10,
         p_wishbone_bd_ram_mem1_197_11, p_wishbone_bd_ram_mem1_197_12,
         p_wishbone_bd_ram_mem1_197_13, p_wishbone_bd_ram_mem1_197_14,
         p_wishbone_bd_ram_mem1_197_15, p_wishbone_bd_ram_mem1_198_8,
         p_wishbone_bd_ram_mem1_198_9, p_wishbone_bd_ram_mem1_198_10,
         p_wishbone_bd_ram_mem1_198_11, p_wishbone_bd_ram_mem1_198_12,
         p_wishbone_bd_ram_mem1_198_13, p_wishbone_bd_ram_mem1_198_14,
         p_wishbone_bd_ram_mem1_198_15, p_wishbone_bd_ram_mem1_199_8,
         p_wishbone_bd_ram_mem1_199_9, p_wishbone_bd_ram_mem1_199_10,
         p_wishbone_bd_ram_mem1_199_11, p_wishbone_bd_ram_mem1_199_12,
         p_wishbone_bd_ram_mem1_199_13, p_wishbone_bd_ram_mem1_199_14,
         p_wishbone_bd_ram_mem1_199_15, p_wishbone_bd_ram_mem1_200_8,
         p_wishbone_bd_ram_mem1_200_9, p_wishbone_bd_ram_mem1_200_10,
         p_wishbone_bd_ram_mem1_200_11, p_wishbone_bd_ram_mem1_200_12,
         p_wishbone_bd_ram_mem1_200_13, p_wishbone_bd_ram_mem1_200_14,
         p_wishbone_bd_ram_mem1_200_15, p_wishbone_bd_ram_mem1_201_8,
         p_wishbone_bd_ram_mem1_201_9, p_wishbone_bd_ram_mem1_201_10,
         p_wishbone_bd_ram_mem1_201_11, p_wishbone_bd_ram_mem1_201_12,
         p_wishbone_bd_ram_mem1_201_13, p_wishbone_bd_ram_mem1_201_14,
         p_wishbone_bd_ram_mem1_201_15, p_wishbone_bd_ram_mem1_202_8,
         p_wishbone_bd_ram_mem1_202_9, p_wishbone_bd_ram_mem1_202_10,
         p_wishbone_bd_ram_mem1_202_11, p_wishbone_bd_ram_mem1_202_12,
         p_wishbone_bd_ram_mem1_202_13, p_wishbone_bd_ram_mem1_202_14,
         p_wishbone_bd_ram_mem1_202_15, p_wishbone_bd_ram_mem1_203_8,
         p_wishbone_bd_ram_mem1_203_9, p_wishbone_bd_ram_mem1_203_10,
         p_wishbone_bd_ram_mem1_203_11, p_wishbone_bd_ram_mem1_203_12,
         p_wishbone_bd_ram_mem1_203_13, p_wishbone_bd_ram_mem1_203_14,
         p_wishbone_bd_ram_mem1_203_15, p_wishbone_bd_ram_mem1_204_8,
         p_wishbone_bd_ram_mem1_204_9, p_wishbone_bd_ram_mem1_204_10,
         p_wishbone_bd_ram_mem1_204_11, p_wishbone_bd_ram_mem1_204_12,
         p_wishbone_bd_ram_mem1_204_13, p_wishbone_bd_ram_mem1_204_14,
         p_wishbone_bd_ram_mem1_204_15, p_wishbone_bd_ram_mem1_205_8,
         p_wishbone_bd_ram_mem1_205_9, p_wishbone_bd_ram_mem1_205_10,
         p_wishbone_bd_ram_mem1_205_11, p_wishbone_bd_ram_mem1_205_12,
         p_wishbone_bd_ram_mem1_205_13, p_wishbone_bd_ram_mem1_205_14,
         p_wishbone_bd_ram_mem1_205_15, p_wishbone_bd_ram_mem1_206_8,
         p_wishbone_bd_ram_mem1_206_9, p_wishbone_bd_ram_mem1_206_10,
         p_wishbone_bd_ram_mem1_206_11, p_wishbone_bd_ram_mem1_206_12,
         p_wishbone_bd_ram_mem1_206_13, p_wishbone_bd_ram_mem1_206_14,
         p_wishbone_bd_ram_mem1_206_15, p_wishbone_bd_ram_mem1_207_8,
         p_wishbone_bd_ram_mem1_207_9, p_wishbone_bd_ram_mem1_207_10,
         p_wishbone_bd_ram_mem1_207_11, p_wishbone_bd_ram_mem1_207_12,
         p_wishbone_bd_ram_mem1_207_13, p_wishbone_bd_ram_mem1_207_14,
         p_wishbone_bd_ram_mem1_207_15, p_wishbone_bd_ram_mem1_208_8,
         p_wishbone_bd_ram_mem1_208_9, p_wishbone_bd_ram_mem1_208_10,
         p_wishbone_bd_ram_mem1_208_11, p_wishbone_bd_ram_mem1_208_12,
         p_wishbone_bd_ram_mem1_208_13, p_wishbone_bd_ram_mem1_208_14,
         p_wishbone_bd_ram_mem1_208_15, p_wishbone_bd_ram_mem1_209_8,
         p_wishbone_bd_ram_mem1_209_9, p_wishbone_bd_ram_mem1_209_10,
         p_wishbone_bd_ram_mem1_209_11, p_wishbone_bd_ram_mem1_209_12,
         p_wishbone_bd_ram_mem1_209_13, p_wishbone_bd_ram_mem1_209_14,
         p_wishbone_bd_ram_mem1_209_15, p_wishbone_bd_ram_mem1_210_8,
         p_wishbone_bd_ram_mem1_210_9, p_wishbone_bd_ram_mem1_210_10,
         p_wishbone_bd_ram_mem1_210_11, p_wishbone_bd_ram_mem1_210_12,
         p_wishbone_bd_ram_mem1_210_13, p_wishbone_bd_ram_mem1_210_14,
         p_wishbone_bd_ram_mem1_210_15, p_wishbone_bd_ram_mem1_211_8,
         p_wishbone_bd_ram_mem1_211_9, p_wishbone_bd_ram_mem1_211_10,
         p_wishbone_bd_ram_mem1_211_11, p_wishbone_bd_ram_mem1_211_12,
         p_wishbone_bd_ram_mem1_211_13, p_wishbone_bd_ram_mem1_211_14,
         p_wishbone_bd_ram_mem1_211_15, p_wishbone_bd_ram_mem1_212_8,
         p_wishbone_bd_ram_mem1_212_9, p_wishbone_bd_ram_mem1_212_10,
         p_wishbone_bd_ram_mem1_212_11, p_wishbone_bd_ram_mem1_212_12,
         p_wishbone_bd_ram_mem1_212_13, p_wishbone_bd_ram_mem1_212_14,
         p_wishbone_bd_ram_mem1_212_15, p_wishbone_bd_ram_mem1_213_8,
         p_wishbone_bd_ram_mem1_213_9, p_wishbone_bd_ram_mem1_213_10,
         p_wishbone_bd_ram_mem1_213_11, p_wishbone_bd_ram_mem1_213_12,
         p_wishbone_bd_ram_mem1_213_13, p_wishbone_bd_ram_mem1_213_14,
         p_wishbone_bd_ram_mem1_213_15, p_wishbone_bd_ram_mem1_214_8,
         p_wishbone_bd_ram_mem1_214_9, p_wishbone_bd_ram_mem1_214_10,
         p_wishbone_bd_ram_mem1_214_11, p_wishbone_bd_ram_mem1_214_12,
         p_wishbone_bd_ram_mem1_214_13, p_wishbone_bd_ram_mem1_214_14,
         p_wishbone_bd_ram_mem1_214_15, p_wishbone_bd_ram_mem1_215_8,
         p_wishbone_bd_ram_mem1_215_9, p_wishbone_bd_ram_mem1_215_10,
         p_wishbone_bd_ram_mem1_215_11, p_wishbone_bd_ram_mem1_215_12,
         p_wishbone_bd_ram_mem1_215_13, p_wishbone_bd_ram_mem1_215_14,
         p_wishbone_bd_ram_mem1_215_15, p_wishbone_bd_ram_mem1_216_8,
         p_wishbone_bd_ram_mem1_216_9, p_wishbone_bd_ram_mem1_216_10,
         p_wishbone_bd_ram_mem1_216_11, p_wishbone_bd_ram_mem1_216_12,
         p_wishbone_bd_ram_mem1_216_13, p_wishbone_bd_ram_mem1_216_14,
         p_wishbone_bd_ram_mem1_216_15, p_wishbone_bd_ram_mem1_217_8,
         p_wishbone_bd_ram_mem1_217_9, p_wishbone_bd_ram_mem1_217_10,
         p_wishbone_bd_ram_mem1_217_11, p_wishbone_bd_ram_mem1_217_12,
         p_wishbone_bd_ram_mem1_217_13, p_wishbone_bd_ram_mem1_217_14,
         p_wishbone_bd_ram_mem1_217_15, p_wishbone_bd_ram_mem1_218_8,
         p_wishbone_bd_ram_mem1_218_9, p_wishbone_bd_ram_mem1_218_10,
         p_wishbone_bd_ram_mem1_218_11, p_wishbone_bd_ram_mem1_218_12,
         p_wishbone_bd_ram_mem1_218_13, p_wishbone_bd_ram_mem1_218_14,
         p_wishbone_bd_ram_mem1_218_15, p_wishbone_bd_ram_mem1_219_8,
         p_wishbone_bd_ram_mem1_219_9, p_wishbone_bd_ram_mem1_219_10,
         p_wishbone_bd_ram_mem1_219_11, p_wishbone_bd_ram_mem1_219_12,
         p_wishbone_bd_ram_mem1_219_13, p_wishbone_bd_ram_mem1_219_14,
         p_wishbone_bd_ram_mem1_219_15, p_wishbone_bd_ram_mem1_220_8,
         p_wishbone_bd_ram_mem1_220_9, p_wishbone_bd_ram_mem1_220_10,
         p_wishbone_bd_ram_mem1_220_11, p_wishbone_bd_ram_mem1_220_12,
         p_wishbone_bd_ram_mem1_220_13, p_wishbone_bd_ram_mem1_220_14,
         p_wishbone_bd_ram_mem1_220_15, p_wishbone_bd_ram_mem1_221_8,
         p_wishbone_bd_ram_mem1_221_9, p_wishbone_bd_ram_mem1_221_10,
         p_wishbone_bd_ram_mem1_221_11, p_wishbone_bd_ram_mem1_221_12,
         p_wishbone_bd_ram_mem1_221_13, p_wishbone_bd_ram_mem1_221_14,
         p_wishbone_bd_ram_mem1_221_15, p_wishbone_bd_ram_mem1_222_8,
         p_wishbone_bd_ram_mem1_222_9, p_wishbone_bd_ram_mem1_222_10,
         p_wishbone_bd_ram_mem1_222_11, p_wishbone_bd_ram_mem1_222_12,
         p_wishbone_bd_ram_mem1_222_13, p_wishbone_bd_ram_mem1_222_14,
         p_wishbone_bd_ram_mem1_222_15, p_wishbone_bd_ram_mem1_223_8,
         p_wishbone_bd_ram_mem1_223_9, p_wishbone_bd_ram_mem1_223_10,
         p_wishbone_bd_ram_mem1_223_11, p_wishbone_bd_ram_mem1_223_12,
         p_wishbone_bd_ram_mem1_223_13, p_wishbone_bd_ram_mem1_223_14,
         p_wishbone_bd_ram_mem1_223_15, p_wishbone_bd_ram_mem1_224_8,
         p_wishbone_bd_ram_mem1_224_9, p_wishbone_bd_ram_mem1_224_10,
         p_wishbone_bd_ram_mem1_224_11, p_wishbone_bd_ram_mem1_224_12,
         p_wishbone_bd_ram_mem1_224_13, p_wishbone_bd_ram_mem1_224_14,
         p_wishbone_bd_ram_mem1_224_15, p_wishbone_bd_ram_mem1_225_8,
         p_wishbone_bd_ram_mem1_225_9, p_wishbone_bd_ram_mem1_225_10,
         p_wishbone_bd_ram_mem1_225_11, p_wishbone_bd_ram_mem1_225_12,
         p_wishbone_bd_ram_mem1_225_13, p_wishbone_bd_ram_mem1_225_14,
         p_wishbone_bd_ram_mem1_225_15, p_wishbone_bd_ram_mem1_226_8,
         p_wishbone_bd_ram_mem1_226_9, p_wishbone_bd_ram_mem1_226_10,
         p_wishbone_bd_ram_mem1_226_11, p_wishbone_bd_ram_mem1_226_12,
         p_wishbone_bd_ram_mem1_226_13, p_wishbone_bd_ram_mem1_226_14,
         p_wishbone_bd_ram_mem1_226_15, p_wishbone_bd_ram_mem1_227_8,
         p_wishbone_bd_ram_mem1_227_9, p_wishbone_bd_ram_mem1_227_10,
         p_wishbone_bd_ram_mem1_227_11, p_wishbone_bd_ram_mem1_227_12,
         p_wishbone_bd_ram_mem1_227_13, p_wishbone_bd_ram_mem1_227_14,
         p_wishbone_bd_ram_mem1_227_15, p_wishbone_bd_ram_mem1_228_8,
         p_wishbone_bd_ram_mem1_228_9, p_wishbone_bd_ram_mem1_228_10,
         p_wishbone_bd_ram_mem1_228_11, p_wishbone_bd_ram_mem1_228_12,
         p_wishbone_bd_ram_mem1_228_13, p_wishbone_bd_ram_mem1_228_14,
         p_wishbone_bd_ram_mem1_228_15, p_wishbone_bd_ram_mem1_229_8,
         p_wishbone_bd_ram_mem1_229_9, p_wishbone_bd_ram_mem1_229_10,
         p_wishbone_bd_ram_mem1_229_11, p_wishbone_bd_ram_mem1_229_12,
         p_wishbone_bd_ram_mem1_229_13, p_wishbone_bd_ram_mem1_229_14,
         p_wishbone_bd_ram_mem1_229_15, p_wishbone_bd_ram_mem1_230_8,
         p_wishbone_bd_ram_mem1_230_9, p_wishbone_bd_ram_mem1_230_10,
         p_wishbone_bd_ram_mem1_230_11, p_wishbone_bd_ram_mem1_230_12,
         p_wishbone_bd_ram_mem1_230_13, p_wishbone_bd_ram_mem1_230_14,
         p_wishbone_bd_ram_mem1_230_15, p_wishbone_bd_ram_mem1_231_8,
         p_wishbone_bd_ram_mem1_231_9, p_wishbone_bd_ram_mem1_231_10,
         p_wishbone_bd_ram_mem1_231_11, p_wishbone_bd_ram_mem1_231_12,
         p_wishbone_bd_ram_mem1_231_13, p_wishbone_bd_ram_mem1_231_14,
         p_wishbone_bd_ram_mem1_231_15, p_wishbone_bd_ram_mem1_232_8,
         p_wishbone_bd_ram_mem1_232_9, p_wishbone_bd_ram_mem1_232_10,
         p_wishbone_bd_ram_mem1_232_11, p_wishbone_bd_ram_mem1_232_12,
         p_wishbone_bd_ram_mem1_232_13, p_wishbone_bd_ram_mem1_232_14,
         p_wishbone_bd_ram_mem1_232_15, p_wishbone_bd_ram_mem1_233_8,
         p_wishbone_bd_ram_mem1_233_9, p_wishbone_bd_ram_mem1_233_10,
         p_wishbone_bd_ram_mem1_233_11, p_wishbone_bd_ram_mem1_233_12,
         p_wishbone_bd_ram_mem1_233_13, p_wishbone_bd_ram_mem1_233_14,
         p_wishbone_bd_ram_mem1_233_15, p_wishbone_bd_ram_mem1_234_8,
         p_wishbone_bd_ram_mem1_234_9, p_wishbone_bd_ram_mem1_234_10,
         p_wishbone_bd_ram_mem1_234_11, p_wishbone_bd_ram_mem1_234_12,
         p_wishbone_bd_ram_mem1_234_13, p_wishbone_bd_ram_mem1_234_14,
         p_wishbone_bd_ram_mem1_234_15, p_wishbone_bd_ram_mem1_235_8,
         p_wishbone_bd_ram_mem1_235_9, p_wishbone_bd_ram_mem1_235_10,
         p_wishbone_bd_ram_mem1_235_11, p_wishbone_bd_ram_mem1_235_12,
         p_wishbone_bd_ram_mem1_235_13, p_wishbone_bd_ram_mem1_235_14,
         p_wishbone_bd_ram_mem1_235_15, p_wishbone_bd_ram_mem1_236_8,
         p_wishbone_bd_ram_mem1_236_9, p_wishbone_bd_ram_mem1_236_10,
         p_wishbone_bd_ram_mem1_236_11, p_wishbone_bd_ram_mem1_236_12,
         p_wishbone_bd_ram_mem1_236_13, p_wishbone_bd_ram_mem1_236_14,
         p_wishbone_bd_ram_mem1_236_15, p_wishbone_bd_ram_mem1_237_8,
         p_wishbone_bd_ram_mem1_237_9, p_wishbone_bd_ram_mem1_237_10,
         p_wishbone_bd_ram_mem1_237_11, p_wishbone_bd_ram_mem1_237_12,
         p_wishbone_bd_ram_mem1_237_13, p_wishbone_bd_ram_mem1_237_14,
         p_wishbone_bd_ram_mem1_237_15, p_wishbone_bd_ram_mem1_238_8,
         p_wishbone_bd_ram_mem1_238_9, p_wishbone_bd_ram_mem1_238_10,
         p_wishbone_bd_ram_mem1_238_11, p_wishbone_bd_ram_mem1_238_12,
         p_wishbone_bd_ram_mem1_238_13, p_wishbone_bd_ram_mem1_238_14,
         p_wishbone_bd_ram_mem1_238_15, p_wishbone_bd_ram_mem1_239_8,
         p_wishbone_bd_ram_mem1_239_9, p_wishbone_bd_ram_mem1_239_10,
         p_wishbone_bd_ram_mem1_239_11, p_wishbone_bd_ram_mem1_239_12,
         p_wishbone_bd_ram_mem1_239_13, p_wishbone_bd_ram_mem1_239_14,
         p_wishbone_bd_ram_mem1_239_15, p_wishbone_bd_ram_mem1_240_8,
         p_wishbone_bd_ram_mem1_240_9, p_wishbone_bd_ram_mem1_240_10,
         p_wishbone_bd_ram_mem1_240_11, p_wishbone_bd_ram_mem1_240_12,
         p_wishbone_bd_ram_mem1_240_13, p_wishbone_bd_ram_mem1_240_14,
         p_wishbone_bd_ram_mem1_240_15, p_wishbone_bd_ram_mem1_241_8,
         p_wishbone_bd_ram_mem1_241_9, p_wishbone_bd_ram_mem1_241_10,
         p_wishbone_bd_ram_mem1_241_11, p_wishbone_bd_ram_mem1_241_12,
         p_wishbone_bd_ram_mem1_241_13, p_wishbone_bd_ram_mem1_241_14,
         p_wishbone_bd_ram_mem1_241_15, p_wishbone_bd_ram_mem1_242_8,
         p_wishbone_bd_ram_mem1_242_9, p_wishbone_bd_ram_mem1_242_10,
         p_wishbone_bd_ram_mem1_242_11, p_wishbone_bd_ram_mem1_242_12,
         p_wishbone_bd_ram_mem1_242_13, p_wishbone_bd_ram_mem1_242_14,
         p_wishbone_bd_ram_mem1_242_15, p_wishbone_bd_ram_mem1_243_8,
         p_wishbone_bd_ram_mem1_243_9, p_wishbone_bd_ram_mem1_243_10,
         p_wishbone_bd_ram_mem1_243_11, p_wishbone_bd_ram_mem1_243_12,
         p_wishbone_bd_ram_mem1_243_13, p_wishbone_bd_ram_mem1_243_14,
         p_wishbone_bd_ram_mem1_243_15, p_wishbone_bd_ram_mem1_244_8,
         p_wishbone_bd_ram_mem1_244_9, p_wishbone_bd_ram_mem1_244_10,
         p_wishbone_bd_ram_mem1_244_11, p_wishbone_bd_ram_mem1_244_12,
         p_wishbone_bd_ram_mem1_244_13, p_wishbone_bd_ram_mem1_244_14,
         p_wishbone_bd_ram_mem1_244_15, p_wishbone_bd_ram_mem1_245_8,
         p_wishbone_bd_ram_mem1_245_9, p_wishbone_bd_ram_mem1_245_10,
         p_wishbone_bd_ram_mem1_245_11, p_wishbone_bd_ram_mem1_245_12,
         p_wishbone_bd_ram_mem1_245_13, p_wishbone_bd_ram_mem1_245_14,
         p_wishbone_bd_ram_mem1_245_15, p_wishbone_bd_ram_mem1_246_8,
         p_wishbone_bd_ram_mem1_246_9, p_wishbone_bd_ram_mem1_246_10,
         p_wishbone_bd_ram_mem1_246_11, p_wishbone_bd_ram_mem1_246_12,
         p_wishbone_bd_ram_mem1_246_13, p_wishbone_bd_ram_mem1_246_14,
         p_wishbone_bd_ram_mem1_246_15, p_wishbone_bd_ram_mem1_247_8,
         p_wishbone_bd_ram_mem1_247_9, p_wishbone_bd_ram_mem1_247_10,
         p_wishbone_bd_ram_mem1_247_11, p_wishbone_bd_ram_mem1_247_12,
         p_wishbone_bd_ram_mem1_247_13, p_wishbone_bd_ram_mem1_247_14,
         p_wishbone_bd_ram_mem1_247_15, p_wishbone_bd_ram_mem1_248_8,
         p_wishbone_bd_ram_mem1_248_9, p_wishbone_bd_ram_mem1_248_10,
         p_wishbone_bd_ram_mem1_248_11, p_wishbone_bd_ram_mem1_248_12,
         p_wishbone_bd_ram_mem1_248_13, p_wishbone_bd_ram_mem1_248_14,
         p_wishbone_bd_ram_mem1_248_15, p_wishbone_bd_ram_mem1_249_8,
         p_wishbone_bd_ram_mem1_249_9, p_wishbone_bd_ram_mem1_249_10,
         p_wishbone_bd_ram_mem1_249_11, p_wishbone_bd_ram_mem1_249_12,
         p_wishbone_bd_ram_mem1_249_13, p_wishbone_bd_ram_mem1_249_14,
         p_wishbone_bd_ram_mem1_249_15, p_wishbone_bd_ram_mem1_250_8,
         p_wishbone_bd_ram_mem1_250_9, p_wishbone_bd_ram_mem1_250_10,
         p_wishbone_bd_ram_mem1_250_11, p_wishbone_bd_ram_mem1_250_12,
         p_wishbone_bd_ram_mem1_250_13, p_wishbone_bd_ram_mem1_250_14,
         p_wishbone_bd_ram_mem1_250_15, p_wishbone_bd_ram_mem1_251_8,
         p_wishbone_bd_ram_mem1_251_9, p_wishbone_bd_ram_mem1_251_10,
         p_wishbone_bd_ram_mem1_251_11, p_wishbone_bd_ram_mem1_251_12,
         p_wishbone_bd_ram_mem1_251_13, p_wishbone_bd_ram_mem1_251_14,
         p_wishbone_bd_ram_mem1_251_15, p_wishbone_bd_ram_mem1_252_8,
         p_wishbone_bd_ram_mem1_252_9, p_wishbone_bd_ram_mem1_252_10,
         p_wishbone_bd_ram_mem1_252_11, p_wishbone_bd_ram_mem1_252_12,
         p_wishbone_bd_ram_mem1_252_13, p_wishbone_bd_ram_mem1_252_14,
         p_wishbone_bd_ram_mem1_252_15, p_wishbone_bd_ram_mem1_253_8,
         p_wishbone_bd_ram_mem1_253_9, p_wishbone_bd_ram_mem1_253_10,
         p_wishbone_bd_ram_mem1_253_11, p_wishbone_bd_ram_mem1_253_12,
         p_wishbone_bd_ram_mem1_253_13, p_wishbone_bd_ram_mem1_253_14,
         p_wishbone_bd_ram_mem1_253_15, p_wishbone_bd_ram_mem1_254_8,
         p_wishbone_bd_ram_mem1_254_9, p_wishbone_bd_ram_mem1_254_10,
         p_wishbone_bd_ram_mem1_254_11, p_wishbone_bd_ram_mem1_254_12,
         p_wishbone_bd_ram_mem1_254_13, p_wishbone_bd_ram_mem1_254_14,
         p_wishbone_bd_ram_mem1_254_15, p_wishbone_bd_ram_mem1_255_8,
         p_wishbone_bd_ram_mem1_255_9, p_wishbone_bd_ram_mem1_255_10,
         p_wishbone_bd_ram_mem1_255_11, p_wishbone_bd_ram_mem1_255_12,
         p_wishbone_bd_ram_mem1_255_13, p_wishbone_bd_ram_mem1_255_14,
         p_wishbone_bd_ram_mem1_255_15, p_wishbone_bd_ram_mem0_0_0,
         p_wishbone_bd_ram_mem0_0_1, p_wishbone_bd_ram_mem0_0_2,
         p_wishbone_bd_ram_mem0_0_3, p_wishbone_bd_ram_mem0_0_4,
         p_wishbone_bd_ram_mem0_0_5, p_wishbone_bd_ram_mem0_0_6,
         p_wishbone_bd_ram_mem0_0_7, p_wishbone_bd_ram_mem0_1_0,
         p_wishbone_bd_ram_mem0_1_1, p_wishbone_bd_ram_mem0_1_2,
         p_wishbone_bd_ram_mem0_1_3, p_wishbone_bd_ram_mem0_1_4,
         p_wishbone_bd_ram_mem0_1_5, p_wishbone_bd_ram_mem0_1_6,
         p_wishbone_bd_ram_mem0_1_7, p_wishbone_bd_ram_mem0_2_0,
         p_wishbone_bd_ram_mem0_2_1, p_wishbone_bd_ram_mem0_2_2,
         p_wishbone_bd_ram_mem0_2_3, p_wishbone_bd_ram_mem0_2_4,
         p_wishbone_bd_ram_mem0_2_5, p_wishbone_bd_ram_mem0_2_6,
         p_wishbone_bd_ram_mem0_2_7, p_wishbone_bd_ram_mem0_3_0,
         p_wishbone_bd_ram_mem0_3_1, p_wishbone_bd_ram_mem0_3_2,
         p_wishbone_bd_ram_mem0_3_3, p_wishbone_bd_ram_mem0_3_4,
         p_wishbone_bd_ram_mem0_3_5, p_wishbone_bd_ram_mem0_3_6,
         p_wishbone_bd_ram_mem0_3_7, p_wishbone_bd_ram_mem0_4_0,
         p_wishbone_bd_ram_mem0_4_1, p_wishbone_bd_ram_mem0_4_2,
         p_wishbone_bd_ram_mem0_4_3, p_wishbone_bd_ram_mem0_4_4,
         p_wishbone_bd_ram_mem0_4_5, p_wishbone_bd_ram_mem0_4_6,
         p_wishbone_bd_ram_mem0_4_7, p_wishbone_bd_ram_mem0_5_0,
         p_wishbone_bd_ram_mem0_5_1, p_wishbone_bd_ram_mem0_5_2,
         p_wishbone_bd_ram_mem0_5_3, p_wishbone_bd_ram_mem0_5_4,
         p_wishbone_bd_ram_mem0_5_5, p_wishbone_bd_ram_mem0_5_6,
         p_wishbone_bd_ram_mem0_5_7, p_wishbone_bd_ram_mem0_6_0,
         p_wishbone_bd_ram_mem0_6_1, p_wishbone_bd_ram_mem0_6_2,
         p_wishbone_bd_ram_mem0_6_3, p_wishbone_bd_ram_mem0_6_4,
         p_wishbone_bd_ram_mem0_6_5, p_wishbone_bd_ram_mem0_6_6,
         p_wishbone_bd_ram_mem0_6_7, p_wishbone_bd_ram_mem0_7_0,
         p_wishbone_bd_ram_mem0_7_1, p_wishbone_bd_ram_mem0_7_2,
         p_wishbone_bd_ram_mem0_7_3, p_wishbone_bd_ram_mem0_7_4,
         p_wishbone_bd_ram_mem0_7_5, p_wishbone_bd_ram_mem0_7_6,
         p_wishbone_bd_ram_mem0_7_7, p_wishbone_bd_ram_mem0_8_0,
         p_wishbone_bd_ram_mem0_8_1, p_wishbone_bd_ram_mem0_8_2,
         p_wishbone_bd_ram_mem0_8_3, p_wishbone_bd_ram_mem0_8_4,
         p_wishbone_bd_ram_mem0_8_5, p_wishbone_bd_ram_mem0_8_6,
         p_wishbone_bd_ram_mem0_8_7, p_wishbone_bd_ram_mem0_9_0,
         p_wishbone_bd_ram_mem0_9_1, p_wishbone_bd_ram_mem0_9_2,
         p_wishbone_bd_ram_mem0_9_3, p_wishbone_bd_ram_mem0_9_4,
         p_wishbone_bd_ram_mem0_9_5, p_wishbone_bd_ram_mem0_9_6,
         p_wishbone_bd_ram_mem0_9_7, p_wishbone_bd_ram_mem0_10_0,
         p_wishbone_bd_ram_mem0_10_1, p_wishbone_bd_ram_mem0_10_2,
         p_wishbone_bd_ram_mem0_10_3, p_wishbone_bd_ram_mem0_10_4,
         p_wishbone_bd_ram_mem0_10_5, p_wishbone_bd_ram_mem0_10_6,
         p_wishbone_bd_ram_mem0_10_7, p_wishbone_bd_ram_mem0_11_0,
         p_wishbone_bd_ram_mem0_11_1, p_wishbone_bd_ram_mem0_11_2,
         p_wishbone_bd_ram_mem0_11_3, p_wishbone_bd_ram_mem0_11_4,
         p_wishbone_bd_ram_mem0_11_5, p_wishbone_bd_ram_mem0_11_6,
         p_wishbone_bd_ram_mem0_11_7, p_wishbone_bd_ram_mem0_12_0,
         p_wishbone_bd_ram_mem0_12_1, p_wishbone_bd_ram_mem0_12_2,
         p_wishbone_bd_ram_mem0_12_3, p_wishbone_bd_ram_mem0_12_4,
         p_wishbone_bd_ram_mem0_12_5, p_wishbone_bd_ram_mem0_12_6,
         p_wishbone_bd_ram_mem0_12_7, p_wishbone_bd_ram_mem0_13_0,
         p_wishbone_bd_ram_mem0_13_1, p_wishbone_bd_ram_mem0_13_2,
         p_wishbone_bd_ram_mem0_13_3, p_wishbone_bd_ram_mem0_13_4,
         p_wishbone_bd_ram_mem0_13_5, p_wishbone_bd_ram_mem0_13_6,
         p_wishbone_bd_ram_mem0_13_7, p_wishbone_bd_ram_mem0_14_0,
         p_wishbone_bd_ram_mem0_14_1, p_wishbone_bd_ram_mem0_14_2,
         p_wishbone_bd_ram_mem0_14_3, p_wishbone_bd_ram_mem0_14_4,
         p_wishbone_bd_ram_mem0_14_5, p_wishbone_bd_ram_mem0_14_6,
         p_wishbone_bd_ram_mem0_14_7, p_wishbone_bd_ram_mem0_15_0,
         p_wishbone_bd_ram_mem0_15_1, p_wishbone_bd_ram_mem0_15_2,
         p_wishbone_bd_ram_mem0_15_3, p_wishbone_bd_ram_mem0_15_4,
         p_wishbone_bd_ram_mem0_15_5, p_wishbone_bd_ram_mem0_15_6,
         p_wishbone_bd_ram_mem0_15_7, p_wishbone_bd_ram_mem0_16_0,
         p_wishbone_bd_ram_mem0_16_1, p_wishbone_bd_ram_mem0_16_2,
         p_wishbone_bd_ram_mem0_16_3, p_wishbone_bd_ram_mem0_16_4,
         p_wishbone_bd_ram_mem0_16_5, p_wishbone_bd_ram_mem0_16_6,
         p_wishbone_bd_ram_mem0_16_7, p_wishbone_bd_ram_mem0_17_0,
         p_wishbone_bd_ram_mem0_17_1, p_wishbone_bd_ram_mem0_17_2,
         p_wishbone_bd_ram_mem0_17_3, p_wishbone_bd_ram_mem0_17_4,
         p_wishbone_bd_ram_mem0_17_5, p_wishbone_bd_ram_mem0_17_6,
         p_wishbone_bd_ram_mem0_17_7, p_wishbone_bd_ram_mem0_18_0,
         p_wishbone_bd_ram_mem0_18_1, p_wishbone_bd_ram_mem0_18_2,
         p_wishbone_bd_ram_mem0_18_3, p_wishbone_bd_ram_mem0_18_4,
         p_wishbone_bd_ram_mem0_18_5, p_wishbone_bd_ram_mem0_18_6,
         p_wishbone_bd_ram_mem0_18_7, p_wishbone_bd_ram_mem0_19_0,
         p_wishbone_bd_ram_mem0_19_1, p_wishbone_bd_ram_mem0_19_2,
         p_wishbone_bd_ram_mem0_19_3, p_wishbone_bd_ram_mem0_19_4,
         p_wishbone_bd_ram_mem0_19_5, p_wishbone_bd_ram_mem0_19_6,
         p_wishbone_bd_ram_mem0_19_7, p_wishbone_bd_ram_mem0_20_0,
         p_wishbone_bd_ram_mem0_20_1, p_wishbone_bd_ram_mem0_20_2,
         p_wishbone_bd_ram_mem0_20_3, p_wishbone_bd_ram_mem0_20_4,
         p_wishbone_bd_ram_mem0_20_5, p_wishbone_bd_ram_mem0_20_6,
         p_wishbone_bd_ram_mem0_20_7, p_wishbone_bd_ram_mem0_21_0,
         p_wishbone_bd_ram_mem0_21_1, p_wishbone_bd_ram_mem0_21_2,
         p_wishbone_bd_ram_mem0_21_3, p_wishbone_bd_ram_mem0_21_4,
         p_wishbone_bd_ram_mem0_21_5, p_wishbone_bd_ram_mem0_21_6,
         p_wishbone_bd_ram_mem0_21_7, p_wishbone_bd_ram_mem0_22_0,
         p_wishbone_bd_ram_mem0_22_1, p_wishbone_bd_ram_mem0_22_2,
         p_wishbone_bd_ram_mem0_22_3, p_wishbone_bd_ram_mem0_22_4,
         p_wishbone_bd_ram_mem0_22_5, p_wishbone_bd_ram_mem0_22_6,
         p_wishbone_bd_ram_mem0_22_7, p_wishbone_bd_ram_mem0_23_0,
         p_wishbone_bd_ram_mem0_23_1, p_wishbone_bd_ram_mem0_23_2,
         p_wishbone_bd_ram_mem0_23_3, p_wishbone_bd_ram_mem0_23_4,
         p_wishbone_bd_ram_mem0_23_5, p_wishbone_bd_ram_mem0_23_6,
         p_wishbone_bd_ram_mem0_23_7, p_wishbone_bd_ram_mem0_24_0,
         p_wishbone_bd_ram_mem0_24_1, p_wishbone_bd_ram_mem0_24_2,
         p_wishbone_bd_ram_mem0_24_3, p_wishbone_bd_ram_mem0_24_4,
         p_wishbone_bd_ram_mem0_24_5, p_wishbone_bd_ram_mem0_24_6,
         p_wishbone_bd_ram_mem0_24_7, p_wishbone_bd_ram_mem0_25_0,
         p_wishbone_bd_ram_mem0_25_1, p_wishbone_bd_ram_mem0_25_2,
         p_wishbone_bd_ram_mem0_25_3, p_wishbone_bd_ram_mem0_25_4,
         p_wishbone_bd_ram_mem0_25_5, p_wishbone_bd_ram_mem0_25_6,
         p_wishbone_bd_ram_mem0_25_7, p_wishbone_bd_ram_mem0_26_0,
         p_wishbone_bd_ram_mem0_26_1, p_wishbone_bd_ram_mem0_26_2,
         p_wishbone_bd_ram_mem0_26_3, p_wishbone_bd_ram_mem0_26_4,
         p_wishbone_bd_ram_mem0_26_5, p_wishbone_bd_ram_mem0_26_6,
         p_wishbone_bd_ram_mem0_26_7, p_wishbone_bd_ram_mem0_27_0,
         p_wishbone_bd_ram_mem0_27_1, p_wishbone_bd_ram_mem0_27_2,
         p_wishbone_bd_ram_mem0_27_3, p_wishbone_bd_ram_mem0_27_4,
         p_wishbone_bd_ram_mem0_27_5, p_wishbone_bd_ram_mem0_27_6,
         p_wishbone_bd_ram_mem0_27_7, p_wishbone_bd_ram_mem0_28_0,
         p_wishbone_bd_ram_mem0_28_1, p_wishbone_bd_ram_mem0_28_2,
         p_wishbone_bd_ram_mem0_28_3, p_wishbone_bd_ram_mem0_28_4,
         p_wishbone_bd_ram_mem0_28_5, p_wishbone_bd_ram_mem0_28_6,
         p_wishbone_bd_ram_mem0_28_7, p_wishbone_bd_ram_mem0_29_0,
         p_wishbone_bd_ram_mem0_29_1, p_wishbone_bd_ram_mem0_29_2,
         p_wishbone_bd_ram_mem0_29_3, p_wishbone_bd_ram_mem0_29_4,
         p_wishbone_bd_ram_mem0_29_5, p_wishbone_bd_ram_mem0_29_6,
         p_wishbone_bd_ram_mem0_29_7, p_wishbone_bd_ram_mem0_30_0,
         p_wishbone_bd_ram_mem0_30_1, p_wishbone_bd_ram_mem0_30_2,
         p_wishbone_bd_ram_mem0_30_3, p_wishbone_bd_ram_mem0_30_4,
         p_wishbone_bd_ram_mem0_30_5, p_wishbone_bd_ram_mem0_30_6,
         p_wishbone_bd_ram_mem0_30_7, p_wishbone_bd_ram_mem0_31_0,
         p_wishbone_bd_ram_mem0_31_1, p_wishbone_bd_ram_mem0_31_2,
         p_wishbone_bd_ram_mem0_31_3, p_wishbone_bd_ram_mem0_31_4,
         p_wishbone_bd_ram_mem0_31_5, p_wishbone_bd_ram_mem0_31_6,
         p_wishbone_bd_ram_mem0_31_7, p_wishbone_bd_ram_mem0_32_0,
         p_wishbone_bd_ram_mem0_32_1, p_wishbone_bd_ram_mem0_32_2,
         p_wishbone_bd_ram_mem0_32_3, p_wishbone_bd_ram_mem0_32_4,
         p_wishbone_bd_ram_mem0_32_5, p_wishbone_bd_ram_mem0_32_6,
         p_wishbone_bd_ram_mem0_32_7, p_wishbone_bd_ram_mem0_33_0,
         p_wishbone_bd_ram_mem0_33_1, p_wishbone_bd_ram_mem0_33_2,
         p_wishbone_bd_ram_mem0_33_3, p_wishbone_bd_ram_mem0_33_4,
         p_wishbone_bd_ram_mem0_33_5, p_wishbone_bd_ram_mem0_33_6,
         p_wishbone_bd_ram_mem0_33_7, p_wishbone_bd_ram_mem0_34_0,
         p_wishbone_bd_ram_mem0_34_1, p_wishbone_bd_ram_mem0_34_2,
         p_wishbone_bd_ram_mem0_34_3, p_wishbone_bd_ram_mem0_34_4,
         p_wishbone_bd_ram_mem0_34_5, p_wishbone_bd_ram_mem0_34_6,
         p_wishbone_bd_ram_mem0_34_7, p_wishbone_bd_ram_mem0_35_0,
         p_wishbone_bd_ram_mem0_35_1, p_wishbone_bd_ram_mem0_35_2,
         p_wishbone_bd_ram_mem0_35_3, p_wishbone_bd_ram_mem0_35_4,
         p_wishbone_bd_ram_mem0_35_5, p_wishbone_bd_ram_mem0_35_6,
         p_wishbone_bd_ram_mem0_35_7, p_wishbone_bd_ram_mem0_36_0,
         p_wishbone_bd_ram_mem0_36_1, p_wishbone_bd_ram_mem0_36_2,
         p_wishbone_bd_ram_mem0_36_3, p_wishbone_bd_ram_mem0_36_4,
         p_wishbone_bd_ram_mem0_36_5, p_wishbone_bd_ram_mem0_36_6,
         p_wishbone_bd_ram_mem0_36_7, p_wishbone_bd_ram_mem0_37_0,
         p_wishbone_bd_ram_mem0_37_1, p_wishbone_bd_ram_mem0_37_2,
         p_wishbone_bd_ram_mem0_37_3, p_wishbone_bd_ram_mem0_37_4,
         p_wishbone_bd_ram_mem0_37_5, p_wishbone_bd_ram_mem0_37_6,
         p_wishbone_bd_ram_mem0_37_7, p_wishbone_bd_ram_mem0_38_0,
         p_wishbone_bd_ram_mem0_38_1, p_wishbone_bd_ram_mem0_38_2,
         p_wishbone_bd_ram_mem0_38_3, p_wishbone_bd_ram_mem0_38_4,
         p_wishbone_bd_ram_mem0_38_5, p_wishbone_bd_ram_mem0_38_6,
         p_wishbone_bd_ram_mem0_38_7, p_wishbone_bd_ram_mem0_39_0,
         p_wishbone_bd_ram_mem0_39_1, p_wishbone_bd_ram_mem0_39_2,
         p_wishbone_bd_ram_mem0_39_3, p_wishbone_bd_ram_mem0_39_4,
         p_wishbone_bd_ram_mem0_39_5, p_wishbone_bd_ram_mem0_39_6,
         p_wishbone_bd_ram_mem0_39_7, p_wishbone_bd_ram_mem0_40_0,
         p_wishbone_bd_ram_mem0_40_1, p_wishbone_bd_ram_mem0_40_2,
         p_wishbone_bd_ram_mem0_40_3, p_wishbone_bd_ram_mem0_40_4,
         p_wishbone_bd_ram_mem0_40_5, p_wishbone_bd_ram_mem0_40_6,
         p_wishbone_bd_ram_mem0_40_7, p_wishbone_bd_ram_mem0_41_0,
         p_wishbone_bd_ram_mem0_41_1, p_wishbone_bd_ram_mem0_41_2,
         p_wishbone_bd_ram_mem0_41_3, p_wishbone_bd_ram_mem0_41_4,
         p_wishbone_bd_ram_mem0_41_5, p_wishbone_bd_ram_mem0_41_6,
         p_wishbone_bd_ram_mem0_41_7, p_wishbone_bd_ram_mem0_42_0,
         p_wishbone_bd_ram_mem0_42_1, p_wishbone_bd_ram_mem0_42_2,
         p_wishbone_bd_ram_mem0_42_3, p_wishbone_bd_ram_mem0_42_4,
         p_wishbone_bd_ram_mem0_42_5, p_wishbone_bd_ram_mem0_42_6,
         p_wishbone_bd_ram_mem0_42_7, p_wishbone_bd_ram_mem0_43_0,
         p_wishbone_bd_ram_mem0_43_1, p_wishbone_bd_ram_mem0_43_2,
         p_wishbone_bd_ram_mem0_43_3, p_wishbone_bd_ram_mem0_43_4,
         p_wishbone_bd_ram_mem0_43_5, p_wishbone_bd_ram_mem0_43_6,
         p_wishbone_bd_ram_mem0_43_7, p_wishbone_bd_ram_mem0_44_0,
         p_wishbone_bd_ram_mem0_44_1, p_wishbone_bd_ram_mem0_44_2,
         p_wishbone_bd_ram_mem0_44_3, p_wishbone_bd_ram_mem0_44_4,
         p_wishbone_bd_ram_mem0_44_5, p_wishbone_bd_ram_mem0_44_6,
         p_wishbone_bd_ram_mem0_44_7, p_wishbone_bd_ram_mem0_45_0,
         p_wishbone_bd_ram_mem0_45_1, p_wishbone_bd_ram_mem0_45_2,
         p_wishbone_bd_ram_mem0_45_3, p_wishbone_bd_ram_mem0_45_4,
         p_wishbone_bd_ram_mem0_45_5, p_wishbone_bd_ram_mem0_45_6,
         p_wishbone_bd_ram_mem0_45_7, p_wishbone_bd_ram_mem0_46_0,
         p_wishbone_bd_ram_mem0_46_1, p_wishbone_bd_ram_mem0_46_2,
         p_wishbone_bd_ram_mem0_46_3, p_wishbone_bd_ram_mem0_46_4,
         p_wishbone_bd_ram_mem0_46_5, p_wishbone_bd_ram_mem0_46_6,
         p_wishbone_bd_ram_mem0_46_7, p_wishbone_bd_ram_mem0_47_0,
         p_wishbone_bd_ram_mem0_47_1, p_wishbone_bd_ram_mem0_47_2,
         p_wishbone_bd_ram_mem0_47_3, p_wishbone_bd_ram_mem0_47_4,
         p_wishbone_bd_ram_mem0_47_5, p_wishbone_bd_ram_mem0_47_6,
         p_wishbone_bd_ram_mem0_47_7, p_wishbone_bd_ram_mem0_48_0,
         p_wishbone_bd_ram_mem0_48_1, p_wishbone_bd_ram_mem0_48_2,
         p_wishbone_bd_ram_mem0_48_3, p_wishbone_bd_ram_mem0_48_4,
         p_wishbone_bd_ram_mem0_48_5, p_wishbone_bd_ram_mem0_48_6,
         p_wishbone_bd_ram_mem0_48_7, p_wishbone_bd_ram_mem0_49_0,
         p_wishbone_bd_ram_mem0_49_1, p_wishbone_bd_ram_mem0_49_2,
         p_wishbone_bd_ram_mem0_49_3, p_wishbone_bd_ram_mem0_49_4,
         p_wishbone_bd_ram_mem0_49_5, p_wishbone_bd_ram_mem0_49_6,
         p_wishbone_bd_ram_mem0_49_7, p_wishbone_bd_ram_mem0_50_0,
         p_wishbone_bd_ram_mem0_50_1, p_wishbone_bd_ram_mem0_50_2,
         p_wishbone_bd_ram_mem0_50_3, p_wishbone_bd_ram_mem0_50_4,
         p_wishbone_bd_ram_mem0_50_5, p_wishbone_bd_ram_mem0_50_6,
         p_wishbone_bd_ram_mem0_50_7, p_wishbone_bd_ram_mem0_51_0,
         p_wishbone_bd_ram_mem0_51_1, p_wishbone_bd_ram_mem0_51_2,
         p_wishbone_bd_ram_mem0_51_3, p_wishbone_bd_ram_mem0_51_4,
         p_wishbone_bd_ram_mem0_51_5, p_wishbone_bd_ram_mem0_51_6,
         p_wishbone_bd_ram_mem0_51_7, p_wishbone_bd_ram_mem0_52_0,
         p_wishbone_bd_ram_mem0_52_1, p_wishbone_bd_ram_mem0_52_2,
         p_wishbone_bd_ram_mem0_52_3, p_wishbone_bd_ram_mem0_52_4,
         p_wishbone_bd_ram_mem0_52_5, p_wishbone_bd_ram_mem0_52_6,
         p_wishbone_bd_ram_mem0_52_7, p_wishbone_bd_ram_mem0_53_0,
         p_wishbone_bd_ram_mem0_53_1, p_wishbone_bd_ram_mem0_53_2,
         p_wishbone_bd_ram_mem0_53_3, p_wishbone_bd_ram_mem0_53_4,
         p_wishbone_bd_ram_mem0_53_5, p_wishbone_bd_ram_mem0_53_6,
         p_wishbone_bd_ram_mem0_53_7, p_wishbone_bd_ram_mem0_54_0,
         p_wishbone_bd_ram_mem0_54_1, p_wishbone_bd_ram_mem0_54_2,
         p_wishbone_bd_ram_mem0_54_3, p_wishbone_bd_ram_mem0_54_4,
         p_wishbone_bd_ram_mem0_54_5, p_wishbone_bd_ram_mem0_54_6,
         p_wishbone_bd_ram_mem0_54_7, p_wishbone_bd_ram_mem0_55_0,
         p_wishbone_bd_ram_mem0_55_1, p_wishbone_bd_ram_mem0_55_2,
         p_wishbone_bd_ram_mem0_55_3, p_wishbone_bd_ram_mem0_55_4,
         p_wishbone_bd_ram_mem0_55_5, p_wishbone_bd_ram_mem0_55_6,
         p_wishbone_bd_ram_mem0_55_7, p_wishbone_bd_ram_mem0_56_0,
         p_wishbone_bd_ram_mem0_56_1, p_wishbone_bd_ram_mem0_56_2,
         p_wishbone_bd_ram_mem0_56_3, p_wishbone_bd_ram_mem0_56_4,
         p_wishbone_bd_ram_mem0_56_5, p_wishbone_bd_ram_mem0_56_6,
         p_wishbone_bd_ram_mem0_56_7, p_wishbone_bd_ram_mem0_57_0,
         p_wishbone_bd_ram_mem0_57_1, p_wishbone_bd_ram_mem0_57_2,
         p_wishbone_bd_ram_mem0_57_3, p_wishbone_bd_ram_mem0_57_4,
         p_wishbone_bd_ram_mem0_57_5, p_wishbone_bd_ram_mem0_57_6,
         p_wishbone_bd_ram_mem0_57_7, p_wishbone_bd_ram_mem0_58_0,
         p_wishbone_bd_ram_mem0_58_1, p_wishbone_bd_ram_mem0_58_2,
         p_wishbone_bd_ram_mem0_58_3, p_wishbone_bd_ram_mem0_58_4,
         p_wishbone_bd_ram_mem0_58_5, p_wishbone_bd_ram_mem0_58_6,
         p_wishbone_bd_ram_mem0_58_7, p_wishbone_bd_ram_mem0_59_0,
         p_wishbone_bd_ram_mem0_59_1, p_wishbone_bd_ram_mem0_59_2,
         p_wishbone_bd_ram_mem0_59_3, p_wishbone_bd_ram_mem0_59_4,
         p_wishbone_bd_ram_mem0_59_5, p_wishbone_bd_ram_mem0_59_6,
         p_wishbone_bd_ram_mem0_59_7, p_wishbone_bd_ram_mem0_60_0,
         p_wishbone_bd_ram_mem0_60_1, p_wishbone_bd_ram_mem0_60_2,
         p_wishbone_bd_ram_mem0_60_3, p_wishbone_bd_ram_mem0_60_4,
         p_wishbone_bd_ram_mem0_60_5, p_wishbone_bd_ram_mem0_60_6,
         p_wishbone_bd_ram_mem0_60_7, p_wishbone_bd_ram_mem0_61_0,
         p_wishbone_bd_ram_mem0_61_1, p_wishbone_bd_ram_mem0_61_2,
         p_wishbone_bd_ram_mem0_61_3, p_wishbone_bd_ram_mem0_61_4,
         p_wishbone_bd_ram_mem0_61_5, p_wishbone_bd_ram_mem0_61_6,
         p_wishbone_bd_ram_mem0_61_7, p_wishbone_bd_ram_mem0_62_0,
         p_wishbone_bd_ram_mem0_62_1, p_wishbone_bd_ram_mem0_62_2,
         p_wishbone_bd_ram_mem0_62_3, p_wishbone_bd_ram_mem0_62_4,
         p_wishbone_bd_ram_mem0_62_5, p_wishbone_bd_ram_mem0_62_6,
         p_wishbone_bd_ram_mem0_62_7, p_wishbone_bd_ram_mem0_63_0,
         p_wishbone_bd_ram_mem0_63_1, p_wishbone_bd_ram_mem0_63_2,
         p_wishbone_bd_ram_mem0_63_3, p_wishbone_bd_ram_mem0_63_4,
         p_wishbone_bd_ram_mem0_63_5, p_wishbone_bd_ram_mem0_63_6,
         p_wishbone_bd_ram_mem0_63_7, p_wishbone_bd_ram_mem0_64_0,
         p_wishbone_bd_ram_mem0_64_1, p_wishbone_bd_ram_mem0_64_2,
         p_wishbone_bd_ram_mem0_64_3, p_wishbone_bd_ram_mem0_64_4,
         p_wishbone_bd_ram_mem0_64_5, p_wishbone_bd_ram_mem0_64_6,
         p_wishbone_bd_ram_mem0_64_7, p_wishbone_bd_ram_mem0_65_0,
         p_wishbone_bd_ram_mem0_65_1, p_wishbone_bd_ram_mem0_65_2,
         p_wishbone_bd_ram_mem0_65_3, p_wishbone_bd_ram_mem0_65_4,
         p_wishbone_bd_ram_mem0_65_5, p_wishbone_bd_ram_mem0_65_6,
         p_wishbone_bd_ram_mem0_65_7, p_wishbone_bd_ram_mem0_66_0,
         p_wishbone_bd_ram_mem0_66_1, p_wishbone_bd_ram_mem0_66_2,
         p_wishbone_bd_ram_mem0_66_3, p_wishbone_bd_ram_mem0_66_4,
         p_wishbone_bd_ram_mem0_66_5, p_wishbone_bd_ram_mem0_66_6,
         p_wishbone_bd_ram_mem0_66_7, p_wishbone_bd_ram_mem0_67_0,
         p_wishbone_bd_ram_mem0_67_1, p_wishbone_bd_ram_mem0_67_2,
         p_wishbone_bd_ram_mem0_67_3, p_wishbone_bd_ram_mem0_67_4,
         p_wishbone_bd_ram_mem0_67_5, p_wishbone_bd_ram_mem0_67_6,
         p_wishbone_bd_ram_mem0_67_7, p_wishbone_bd_ram_mem0_68_0,
         p_wishbone_bd_ram_mem0_68_1, p_wishbone_bd_ram_mem0_68_2,
         p_wishbone_bd_ram_mem0_68_3, p_wishbone_bd_ram_mem0_68_4,
         p_wishbone_bd_ram_mem0_68_5, p_wishbone_bd_ram_mem0_68_6,
         p_wishbone_bd_ram_mem0_68_7, p_wishbone_bd_ram_mem0_69_0,
         p_wishbone_bd_ram_mem0_69_1, p_wishbone_bd_ram_mem0_69_2,
         p_wishbone_bd_ram_mem0_69_3, p_wishbone_bd_ram_mem0_69_4,
         p_wishbone_bd_ram_mem0_69_5, p_wishbone_bd_ram_mem0_69_6,
         p_wishbone_bd_ram_mem0_69_7, p_wishbone_bd_ram_mem0_70_0,
         p_wishbone_bd_ram_mem0_70_1, p_wishbone_bd_ram_mem0_70_2,
         p_wishbone_bd_ram_mem0_70_3, p_wishbone_bd_ram_mem0_70_4,
         p_wishbone_bd_ram_mem0_70_5, p_wishbone_bd_ram_mem0_70_6,
         p_wishbone_bd_ram_mem0_70_7, p_wishbone_bd_ram_mem0_71_0,
         p_wishbone_bd_ram_mem0_71_1, p_wishbone_bd_ram_mem0_71_2,
         p_wishbone_bd_ram_mem0_71_3, p_wishbone_bd_ram_mem0_71_4,
         p_wishbone_bd_ram_mem0_71_5, p_wishbone_bd_ram_mem0_71_6,
         p_wishbone_bd_ram_mem0_71_7, p_wishbone_bd_ram_mem0_72_0,
         p_wishbone_bd_ram_mem0_72_1, p_wishbone_bd_ram_mem0_72_2,
         p_wishbone_bd_ram_mem0_72_3, p_wishbone_bd_ram_mem0_72_4,
         p_wishbone_bd_ram_mem0_72_5, p_wishbone_bd_ram_mem0_72_6,
         p_wishbone_bd_ram_mem0_72_7, p_wishbone_bd_ram_mem0_73_0,
         p_wishbone_bd_ram_mem0_73_1, p_wishbone_bd_ram_mem0_73_2,
         p_wishbone_bd_ram_mem0_73_3, p_wishbone_bd_ram_mem0_73_4,
         p_wishbone_bd_ram_mem0_73_5, p_wishbone_bd_ram_mem0_73_6,
         p_wishbone_bd_ram_mem0_73_7, p_wishbone_bd_ram_mem0_74_0,
         p_wishbone_bd_ram_mem0_74_1, p_wishbone_bd_ram_mem0_74_2,
         p_wishbone_bd_ram_mem0_74_3, p_wishbone_bd_ram_mem0_74_4,
         p_wishbone_bd_ram_mem0_74_5, p_wishbone_bd_ram_mem0_74_6,
         p_wishbone_bd_ram_mem0_74_7, p_wishbone_bd_ram_mem0_75_0,
         p_wishbone_bd_ram_mem0_75_1, p_wishbone_bd_ram_mem0_75_2,
         p_wishbone_bd_ram_mem0_75_3, p_wishbone_bd_ram_mem0_75_4,
         p_wishbone_bd_ram_mem0_75_5, p_wishbone_bd_ram_mem0_75_6,
         p_wishbone_bd_ram_mem0_75_7, p_wishbone_bd_ram_mem0_76_0,
         p_wishbone_bd_ram_mem0_76_1, p_wishbone_bd_ram_mem0_76_2,
         p_wishbone_bd_ram_mem0_76_3, p_wishbone_bd_ram_mem0_76_4,
         p_wishbone_bd_ram_mem0_76_5, p_wishbone_bd_ram_mem0_76_6,
         p_wishbone_bd_ram_mem0_76_7, p_wishbone_bd_ram_mem0_77_0,
         p_wishbone_bd_ram_mem0_77_1, p_wishbone_bd_ram_mem0_77_2,
         p_wishbone_bd_ram_mem0_77_3, p_wishbone_bd_ram_mem0_77_4,
         p_wishbone_bd_ram_mem0_77_5, p_wishbone_bd_ram_mem0_77_6,
         p_wishbone_bd_ram_mem0_77_7, p_wishbone_bd_ram_mem0_78_0,
         p_wishbone_bd_ram_mem0_78_1, p_wishbone_bd_ram_mem0_78_2,
         p_wishbone_bd_ram_mem0_78_3, p_wishbone_bd_ram_mem0_78_4,
         p_wishbone_bd_ram_mem0_78_5, p_wishbone_bd_ram_mem0_78_6,
         p_wishbone_bd_ram_mem0_78_7, p_wishbone_bd_ram_mem0_79_0,
         p_wishbone_bd_ram_mem0_79_1, p_wishbone_bd_ram_mem0_79_2,
         p_wishbone_bd_ram_mem0_79_3, p_wishbone_bd_ram_mem0_79_4,
         p_wishbone_bd_ram_mem0_79_5, p_wishbone_bd_ram_mem0_79_6,
         p_wishbone_bd_ram_mem0_79_7, p_wishbone_bd_ram_mem0_80_0,
         p_wishbone_bd_ram_mem0_80_1, p_wishbone_bd_ram_mem0_80_2,
         p_wishbone_bd_ram_mem0_80_3, p_wishbone_bd_ram_mem0_80_4,
         p_wishbone_bd_ram_mem0_80_5, p_wishbone_bd_ram_mem0_80_6,
         p_wishbone_bd_ram_mem0_80_7, p_wishbone_bd_ram_mem0_81_0,
         p_wishbone_bd_ram_mem0_81_1, p_wishbone_bd_ram_mem0_81_2,
         p_wishbone_bd_ram_mem0_81_3, p_wishbone_bd_ram_mem0_81_4,
         p_wishbone_bd_ram_mem0_81_5, p_wishbone_bd_ram_mem0_81_6,
         p_wishbone_bd_ram_mem0_81_7, p_wishbone_bd_ram_mem0_82_0,
         p_wishbone_bd_ram_mem0_82_1, p_wishbone_bd_ram_mem0_82_2,
         p_wishbone_bd_ram_mem0_82_3, p_wishbone_bd_ram_mem0_82_4,
         p_wishbone_bd_ram_mem0_82_5, p_wishbone_bd_ram_mem0_82_6,
         p_wishbone_bd_ram_mem0_82_7, p_wishbone_bd_ram_mem0_83_0,
         p_wishbone_bd_ram_mem0_83_1, p_wishbone_bd_ram_mem0_83_2,
         p_wishbone_bd_ram_mem0_83_3, p_wishbone_bd_ram_mem0_83_4,
         p_wishbone_bd_ram_mem0_83_5, p_wishbone_bd_ram_mem0_83_6,
         p_wishbone_bd_ram_mem0_83_7, p_wishbone_bd_ram_mem0_84_0,
         p_wishbone_bd_ram_mem0_84_1, p_wishbone_bd_ram_mem0_84_2,
         p_wishbone_bd_ram_mem0_84_3, p_wishbone_bd_ram_mem0_84_4,
         p_wishbone_bd_ram_mem0_84_5, p_wishbone_bd_ram_mem0_84_6,
         p_wishbone_bd_ram_mem0_84_7, p_wishbone_bd_ram_mem0_85_0,
         p_wishbone_bd_ram_mem0_85_1, p_wishbone_bd_ram_mem0_85_2,
         p_wishbone_bd_ram_mem0_85_3, p_wishbone_bd_ram_mem0_85_4,
         p_wishbone_bd_ram_mem0_85_5, p_wishbone_bd_ram_mem0_85_6,
         p_wishbone_bd_ram_mem0_85_7, p_wishbone_bd_ram_mem0_86_0,
         p_wishbone_bd_ram_mem0_86_1, p_wishbone_bd_ram_mem0_86_2,
         p_wishbone_bd_ram_mem0_86_3, p_wishbone_bd_ram_mem0_86_4,
         p_wishbone_bd_ram_mem0_86_5, p_wishbone_bd_ram_mem0_86_6,
         p_wishbone_bd_ram_mem0_86_7, p_wishbone_bd_ram_mem0_87_0,
         p_wishbone_bd_ram_mem0_87_1, p_wishbone_bd_ram_mem0_87_2,
         p_wishbone_bd_ram_mem0_87_3, p_wishbone_bd_ram_mem0_87_4,
         p_wishbone_bd_ram_mem0_87_5, p_wishbone_bd_ram_mem0_87_6,
         p_wishbone_bd_ram_mem0_87_7, p_wishbone_bd_ram_mem0_88_0,
         p_wishbone_bd_ram_mem0_88_1, p_wishbone_bd_ram_mem0_88_2,
         p_wishbone_bd_ram_mem0_88_3, p_wishbone_bd_ram_mem0_88_4,
         p_wishbone_bd_ram_mem0_88_5, p_wishbone_bd_ram_mem0_88_6,
         p_wishbone_bd_ram_mem0_88_7, p_wishbone_bd_ram_mem0_89_0,
         p_wishbone_bd_ram_mem0_89_1, p_wishbone_bd_ram_mem0_89_2,
         p_wishbone_bd_ram_mem0_89_3, p_wishbone_bd_ram_mem0_89_4,
         p_wishbone_bd_ram_mem0_89_5, p_wishbone_bd_ram_mem0_89_6,
         p_wishbone_bd_ram_mem0_89_7, p_wishbone_bd_ram_mem0_90_0,
         p_wishbone_bd_ram_mem0_90_1, p_wishbone_bd_ram_mem0_90_2,
         p_wishbone_bd_ram_mem0_90_3, p_wishbone_bd_ram_mem0_90_4,
         p_wishbone_bd_ram_mem0_90_5, p_wishbone_bd_ram_mem0_90_6,
         p_wishbone_bd_ram_mem0_90_7, p_wishbone_bd_ram_mem0_91_0,
         p_wishbone_bd_ram_mem0_91_1, p_wishbone_bd_ram_mem0_91_2,
         p_wishbone_bd_ram_mem0_91_3, p_wishbone_bd_ram_mem0_91_4,
         p_wishbone_bd_ram_mem0_91_5, p_wishbone_bd_ram_mem0_91_6,
         p_wishbone_bd_ram_mem0_91_7, p_wishbone_bd_ram_mem0_92_0,
         p_wishbone_bd_ram_mem0_92_1, p_wishbone_bd_ram_mem0_92_2,
         p_wishbone_bd_ram_mem0_92_3, p_wishbone_bd_ram_mem0_92_4,
         p_wishbone_bd_ram_mem0_92_5, p_wishbone_bd_ram_mem0_92_6,
         p_wishbone_bd_ram_mem0_92_7, p_wishbone_bd_ram_mem0_93_0,
         p_wishbone_bd_ram_mem0_93_1, p_wishbone_bd_ram_mem0_93_2,
         p_wishbone_bd_ram_mem0_93_3, p_wishbone_bd_ram_mem0_93_4,
         p_wishbone_bd_ram_mem0_93_5, p_wishbone_bd_ram_mem0_93_6,
         p_wishbone_bd_ram_mem0_93_7, p_wishbone_bd_ram_mem0_94_0,
         p_wishbone_bd_ram_mem0_94_1, p_wishbone_bd_ram_mem0_94_2,
         p_wishbone_bd_ram_mem0_94_3, p_wishbone_bd_ram_mem0_94_4,
         p_wishbone_bd_ram_mem0_94_5, p_wishbone_bd_ram_mem0_94_6,
         p_wishbone_bd_ram_mem0_94_7, p_wishbone_bd_ram_mem0_95_0,
         p_wishbone_bd_ram_mem0_95_1, p_wishbone_bd_ram_mem0_95_2,
         p_wishbone_bd_ram_mem0_95_3, p_wishbone_bd_ram_mem0_95_4,
         p_wishbone_bd_ram_mem0_95_5, p_wishbone_bd_ram_mem0_95_6,
         p_wishbone_bd_ram_mem0_95_7, p_wishbone_bd_ram_mem0_96_0,
         p_wishbone_bd_ram_mem0_96_1, p_wishbone_bd_ram_mem0_96_2,
         p_wishbone_bd_ram_mem0_96_3, p_wishbone_bd_ram_mem0_96_4,
         p_wishbone_bd_ram_mem0_96_5, p_wishbone_bd_ram_mem0_96_6,
         p_wishbone_bd_ram_mem0_96_7, p_wishbone_bd_ram_mem0_97_0,
         p_wishbone_bd_ram_mem0_97_1, p_wishbone_bd_ram_mem0_97_2,
         p_wishbone_bd_ram_mem0_97_3, p_wishbone_bd_ram_mem0_97_4,
         p_wishbone_bd_ram_mem0_97_5, p_wishbone_bd_ram_mem0_97_6,
         p_wishbone_bd_ram_mem0_97_7, p_wishbone_bd_ram_mem0_98_0,
         p_wishbone_bd_ram_mem0_98_1, p_wishbone_bd_ram_mem0_98_2,
         p_wishbone_bd_ram_mem0_98_3, p_wishbone_bd_ram_mem0_98_4,
         p_wishbone_bd_ram_mem0_98_5, p_wishbone_bd_ram_mem0_98_6,
         p_wishbone_bd_ram_mem0_98_7, p_wishbone_bd_ram_mem0_99_0,
         p_wishbone_bd_ram_mem0_99_1, p_wishbone_bd_ram_mem0_99_2,
         p_wishbone_bd_ram_mem0_99_3, p_wishbone_bd_ram_mem0_99_4,
         p_wishbone_bd_ram_mem0_99_5, p_wishbone_bd_ram_mem0_99_6,
         p_wishbone_bd_ram_mem0_99_7, p_wishbone_bd_ram_mem0_100_0,
         p_wishbone_bd_ram_mem0_100_1, p_wishbone_bd_ram_mem0_100_2,
         p_wishbone_bd_ram_mem0_100_3, p_wishbone_bd_ram_mem0_100_4,
         p_wishbone_bd_ram_mem0_100_5, p_wishbone_bd_ram_mem0_100_6,
         p_wishbone_bd_ram_mem0_100_7, p_wishbone_bd_ram_mem0_101_0,
         p_wishbone_bd_ram_mem0_101_1, p_wishbone_bd_ram_mem0_101_2,
         p_wishbone_bd_ram_mem0_101_3, p_wishbone_bd_ram_mem0_101_4,
         p_wishbone_bd_ram_mem0_101_5, p_wishbone_bd_ram_mem0_101_6,
         p_wishbone_bd_ram_mem0_101_7, p_wishbone_bd_ram_mem0_102_0,
         p_wishbone_bd_ram_mem0_102_1, p_wishbone_bd_ram_mem0_102_2,
         p_wishbone_bd_ram_mem0_102_3, p_wishbone_bd_ram_mem0_102_4,
         p_wishbone_bd_ram_mem0_102_5, p_wishbone_bd_ram_mem0_102_6,
         p_wishbone_bd_ram_mem0_102_7, p_wishbone_bd_ram_mem0_103_0,
         p_wishbone_bd_ram_mem0_103_1, p_wishbone_bd_ram_mem0_103_2,
         p_wishbone_bd_ram_mem0_103_3, p_wishbone_bd_ram_mem0_103_4,
         p_wishbone_bd_ram_mem0_103_5, p_wishbone_bd_ram_mem0_103_6,
         p_wishbone_bd_ram_mem0_103_7, p_wishbone_bd_ram_mem0_104_0,
         p_wishbone_bd_ram_mem0_104_1, p_wishbone_bd_ram_mem0_104_2,
         p_wishbone_bd_ram_mem0_104_3, p_wishbone_bd_ram_mem0_104_4,
         p_wishbone_bd_ram_mem0_104_5, p_wishbone_bd_ram_mem0_104_6,
         p_wishbone_bd_ram_mem0_104_7, p_wishbone_bd_ram_mem0_105_0,
         p_wishbone_bd_ram_mem0_105_1, p_wishbone_bd_ram_mem0_105_2,
         p_wishbone_bd_ram_mem0_105_3, p_wishbone_bd_ram_mem0_105_4,
         p_wishbone_bd_ram_mem0_105_5, p_wishbone_bd_ram_mem0_105_6,
         p_wishbone_bd_ram_mem0_105_7, p_wishbone_bd_ram_mem0_106_0,
         p_wishbone_bd_ram_mem0_106_1, p_wishbone_bd_ram_mem0_106_2,
         p_wishbone_bd_ram_mem0_106_3, p_wishbone_bd_ram_mem0_106_4,
         p_wishbone_bd_ram_mem0_106_5, p_wishbone_bd_ram_mem0_106_6,
         p_wishbone_bd_ram_mem0_106_7, p_wishbone_bd_ram_mem0_107_0,
         p_wishbone_bd_ram_mem0_107_1, p_wishbone_bd_ram_mem0_107_2,
         p_wishbone_bd_ram_mem0_107_3, p_wishbone_bd_ram_mem0_107_4,
         p_wishbone_bd_ram_mem0_107_5, p_wishbone_bd_ram_mem0_107_6,
         p_wishbone_bd_ram_mem0_107_7, p_wishbone_bd_ram_mem0_108_0,
         p_wishbone_bd_ram_mem0_108_1, p_wishbone_bd_ram_mem0_108_2,
         p_wishbone_bd_ram_mem0_108_3, p_wishbone_bd_ram_mem0_108_4,
         p_wishbone_bd_ram_mem0_108_5, p_wishbone_bd_ram_mem0_108_6,
         p_wishbone_bd_ram_mem0_108_7, p_wishbone_bd_ram_mem0_109_0,
         p_wishbone_bd_ram_mem0_109_1, p_wishbone_bd_ram_mem0_109_2,
         p_wishbone_bd_ram_mem0_109_3, p_wishbone_bd_ram_mem0_109_4,
         p_wishbone_bd_ram_mem0_109_5, p_wishbone_bd_ram_mem0_109_6,
         p_wishbone_bd_ram_mem0_109_7, p_wishbone_bd_ram_mem0_110_0,
         p_wishbone_bd_ram_mem0_110_1, p_wishbone_bd_ram_mem0_110_2,
         p_wishbone_bd_ram_mem0_110_3, p_wishbone_bd_ram_mem0_110_4,
         p_wishbone_bd_ram_mem0_110_5, p_wishbone_bd_ram_mem0_110_6,
         p_wishbone_bd_ram_mem0_110_7, p_wishbone_bd_ram_mem0_111_0,
         p_wishbone_bd_ram_mem0_111_1, p_wishbone_bd_ram_mem0_111_2,
         p_wishbone_bd_ram_mem0_111_3, p_wishbone_bd_ram_mem0_111_4,
         p_wishbone_bd_ram_mem0_111_5, p_wishbone_bd_ram_mem0_111_6,
         p_wishbone_bd_ram_mem0_111_7, p_wishbone_bd_ram_mem0_112_0,
         p_wishbone_bd_ram_mem0_112_1, p_wishbone_bd_ram_mem0_112_2,
         p_wishbone_bd_ram_mem0_112_3, p_wishbone_bd_ram_mem0_112_4,
         p_wishbone_bd_ram_mem0_112_5, p_wishbone_bd_ram_mem0_112_6,
         p_wishbone_bd_ram_mem0_112_7, p_wishbone_bd_ram_mem0_113_0,
         p_wishbone_bd_ram_mem0_113_1, p_wishbone_bd_ram_mem0_113_2,
         p_wishbone_bd_ram_mem0_113_3, p_wishbone_bd_ram_mem0_113_4,
         p_wishbone_bd_ram_mem0_113_5, p_wishbone_bd_ram_mem0_113_6,
         p_wishbone_bd_ram_mem0_113_7, p_wishbone_bd_ram_mem0_114_0,
         p_wishbone_bd_ram_mem0_114_1, p_wishbone_bd_ram_mem0_114_2,
         p_wishbone_bd_ram_mem0_114_3, p_wishbone_bd_ram_mem0_114_4,
         p_wishbone_bd_ram_mem0_114_5, p_wishbone_bd_ram_mem0_114_6,
         p_wishbone_bd_ram_mem0_114_7, p_wishbone_bd_ram_mem0_115_0,
         p_wishbone_bd_ram_mem0_115_1, p_wishbone_bd_ram_mem0_115_2,
         p_wishbone_bd_ram_mem0_115_3, p_wishbone_bd_ram_mem0_115_4,
         p_wishbone_bd_ram_mem0_115_5, p_wishbone_bd_ram_mem0_115_6,
         p_wishbone_bd_ram_mem0_115_7, p_wishbone_bd_ram_mem0_116_0,
         p_wishbone_bd_ram_mem0_116_1, p_wishbone_bd_ram_mem0_116_2,
         p_wishbone_bd_ram_mem0_116_3, p_wishbone_bd_ram_mem0_116_4,
         p_wishbone_bd_ram_mem0_116_5, p_wishbone_bd_ram_mem0_116_6,
         p_wishbone_bd_ram_mem0_116_7, p_wishbone_bd_ram_mem0_117_0,
         p_wishbone_bd_ram_mem0_117_1, p_wishbone_bd_ram_mem0_117_2,
         p_wishbone_bd_ram_mem0_117_3, p_wishbone_bd_ram_mem0_117_4,
         p_wishbone_bd_ram_mem0_117_5, p_wishbone_bd_ram_mem0_117_6,
         p_wishbone_bd_ram_mem0_117_7, p_wishbone_bd_ram_mem0_118_0,
         p_wishbone_bd_ram_mem0_118_1, p_wishbone_bd_ram_mem0_118_2,
         p_wishbone_bd_ram_mem0_118_3, p_wishbone_bd_ram_mem0_118_4,
         p_wishbone_bd_ram_mem0_118_5, p_wishbone_bd_ram_mem0_118_6,
         p_wishbone_bd_ram_mem0_118_7, p_wishbone_bd_ram_mem0_119_0,
         p_wishbone_bd_ram_mem0_119_1, p_wishbone_bd_ram_mem0_119_2,
         p_wishbone_bd_ram_mem0_119_3, p_wishbone_bd_ram_mem0_119_4,
         p_wishbone_bd_ram_mem0_119_5, p_wishbone_bd_ram_mem0_119_6,
         p_wishbone_bd_ram_mem0_119_7, p_wishbone_bd_ram_mem0_120_0,
         p_wishbone_bd_ram_mem0_120_1, p_wishbone_bd_ram_mem0_120_2,
         p_wishbone_bd_ram_mem0_120_3, p_wishbone_bd_ram_mem0_120_4,
         p_wishbone_bd_ram_mem0_120_5, p_wishbone_bd_ram_mem0_120_6,
         p_wishbone_bd_ram_mem0_120_7, p_wishbone_bd_ram_mem0_121_0,
         p_wishbone_bd_ram_mem0_121_1, p_wishbone_bd_ram_mem0_121_2,
         p_wishbone_bd_ram_mem0_121_3, p_wishbone_bd_ram_mem0_121_4,
         p_wishbone_bd_ram_mem0_121_5, p_wishbone_bd_ram_mem0_121_6,
         p_wishbone_bd_ram_mem0_121_7, p_wishbone_bd_ram_mem0_122_0,
         p_wishbone_bd_ram_mem0_122_1, p_wishbone_bd_ram_mem0_122_2,
         p_wishbone_bd_ram_mem0_122_3, p_wishbone_bd_ram_mem0_122_4,
         p_wishbone_bd_ram_mem0_122_5, p_wishbone_bd_ram_mem0_122_6,
         p_wishbone_bd_ram_mem0_122_7, p_wishbone_bd_ram_mem0_123_0,
         p_wishbone_bd_ram_mem0_123_1, p_wishbone_bd_ram_mem0_123_2,
         p_wishbone_bd_ram_mem0_123_3, p_wishbone_bd_ram_mem0_123_4,
         p_wishbone_bd_ram_mem0_123_5, p_wishbone_bd_ram_mem0_123_6,
         p_wishbone_bd_ram_mem0_123_7, p_wishbone_bd_ram_mem0_124_0,
         p_wishbone_bd_ram_mem0_124_1, p_wishbone_bd_ram_mem0_124_2,
         p_wishbone_bd_ram_mem0_124_3, p_wishbone_bd_ram_mem0_124_4,
         p_wishbone_bd_ram_mem0_124_5, p_wishbone_bd_ram_mem0_124_6,
         p_wishbone_bd_ram_mem0_124_7, p_wishbone_bd_ram_mem0_125_0,
         p_wishbone_bd_ram_mem0_125_1, p_wishbone_bd_ram_mem0_125_2,
         p_wishbone_bd_ram_mem0_125_3, p_wishbone_bd_ram_mem0_125_4,
         p_wishbone_bd_ram_mem0_125_5, p_wishbone_bd_ram_mem0_125_6,
         p_wishbone_bd_ram_mem0_125_7, p_wishbone_bd_ram_mem0_126_0,
         p_wishbone_bd_ram_mem0_126_1, p_wishbone_bd_ram_mem0_126_2,
         p_wishbone_bd_ram_mem0_126_3, p_wishbone_bd_ram_mem0_126_4,
         p_wishbone_bd_ram_mem0_126_5, p_wishbone_bd_ram_mem0_126_6,
         p_wishbone_bd_ram_mem0_126_7, p_wishbone_bd_ram_mem0_127_0,
         p_wishbone_bd_ram_mem0_127_1, p_wishbone_bd_ram_mem0_127_2,
         p_wishbone_bd_ram_mem0_127_3, p_wishbone_bd_ram_mem0_127_4,
         p_wishbone_bd_ram_mem0_127_5, p_wishbone_bd_ram_mem0_127_6,
         p_wishbone_bd_ram_mem0_127_7, p_wishbone_bd_ram_mem0_128_0,
         p_wishbone_bd_ram_mem0_128_1, p_wishbone_bd_ram_mem0_128_2,
         p_wishbone_bd_ram_mem0_128_3, p_wishbone_bd_ram_mem0_128_4,
         p_wishbone_bd_ram_mem0_128_5, p_wishbone_bd_ram_mem0_128_6,
         p_wishbone_bd_ram_mem0_128_7, p_wishbone_bd_ram_mem0_129_0,
         p_wishbone_bd_ram_mem0_129_1, p_wishbone_bd_ram_mem0_129_2,
         p_wishbone_bd_ram_mem0_129_3, p_wishbone_bd_ram_mem0_129_4,
         p_wishbone_bd_ram_mem0_129_5, p_wishbone_bd_ram_mem0_129_6,
         p_wishbone_bd_ram_mem0_129_7, p_wishbone_bd_ram_mem0_130_0,
         p_wishbone_bd_ram_mem0_130_1, p_wishbone_bd_ram_mem0_130_2,
         p_wishbone_bd_ram_mem0_130_3, p_wishbone_bd_ram_mem0_130_4,
         p_wishbone_bd_ram_mem0_130_5, p_wishbone_bd_ram_mem0_130_6,
         p_wishbone_bd_ram_mem0_130_7, p_wishbone_bd_ram_mem0_131_0,
         p_wishbone_bd_ram_mem0_131_1, p_wishbone_bd_ram_mem0_131_2,
         p_wishbone_bd_ram_mem0_131_3, p_wishbone_bd_ram_mem0_131_4,
         p_wishbone_bd_ram_mem0_131_5, p_wishbone_bd_ram_mem0_131_6,
         p_wishbone_bd_ram_mem0_131_7, p_wishbone_bd_ram_mem0_132_0,
         p_wishbone_bd_ram_mem0_132_1, p_wishbone_bd_ram_mem0_132_2,
         p_wishbone_bd_ram_mem0_132_3, p_wishbone_bd_ram_mem0_132_4,
         p_wishbone_bd_ram_mem0_132_5, p_wishbone_bd_ram_mem0_132_6,
         p_wishbone_bd_ram_mem0_132_7, p_wishbone_bd_ram_mem0_133_0,
         p_wishbone_bd_ram_mem0_133_1, p_wishbone_bd_ram_mem0_133_2,
         p_wishbone_bd_ram_mem0_133_3, p_wishbone_bd_ram_mem0_133_4,
         p_wishbone_bd_ram_mem0_133_5, p_wishbone_bd_ram_mem0_133_6,
         p_wishbone_bd_ram_mem0_133_7, p_wishbone_bd_ram_mem0_134_0,
         p_wishbone_bd_ram_mem0_134_1, p_wishbone_bd_ram_mem0_134_2,
         p_wishbone_bd_ram_mem0_134_3, p_wishbone_bd_ram_mem0_134_4,
         p_wishbone_bd_ram_mem0_134_5, p_wishbone_bd_ram_mem0_134_6,
         p_wishbone_bd_ram_mem0_134_7, p_wishbone_bd_ram_mem0_135_0,
         p_wishbone_bd_ram_mem0_135_1, p_wishbone_bd_ram_mem0_135_2,
         p_wishbone_bd_ram_mem0_135_3, p_wishbone_bd_ram_mem0_135_4,
         p_wishbone_bd_ram_mem0_135_5, p_wishbone_bd_ram_mem0_135_6,
         p_wishbone_bd_ram_mem0_135_7, p_wishbone_bd_ram_mem0_136_0,
         p_wishbone_bd_ram_mem0_136_1, p_wishbone_bd_ram_mem0_136_2,
         p_wishbone_bd_ram_mem0_136_3, p_wishbone_bd_ram_mem0_136_4,
         p_wishbone_bd_ram_mem0_136_5, p_wishbone_bd_ram_mem0_136_6,
         p_wishbone_bd_ram_mem0_136_7, p_wishbone_bd_ram_mem0_137_0,
         p_wishbone_bd_ram_mem0_137_1, p_wishbone_bd_ram_mem0_137_2,
         p_wishbone_bd_ram_mem0_137_3, p_wishbone_bd_ram_mem0_137_4,
         p_wishbone_bd_ram_mem0_137_5, p_wishbone_bd_ram_mem0_137_6,
         p_wishbone_bd_ram_mem0_137_7, p_wishbone_bd_ram_mem0_138_0,
         p_wishbone_bd_ram_mem0_138_1, p_wishbone_bd_ram_mem0_138_2,
         p_wishbone_bd_ram_mem0_138_3, p_wishbone_bd_ram_mem0_138_4,
         p_wishbone_bd_ram_mem0_138_5, p_wishbone_bd_ram_mem0_138_6,
         p_wishbone_bd_ram_mem0_138_7, p_wishbone_bd_ram_mem0_139_0,
         p_wishbone_bd_ram_mem0_139_1, p_wishbone_bd_ram_mem0_139_2,
         p_wishbone_bd_ram_mem0_139_3, p_wishbone_bd_ram_mem0_139_4,
         p_wishbone_bd_ram_mem0_139_5, p_wishbone_bd_ram_mem0_139_6,
         p_wishbone_bd_ram_mem0_139_7, p_wishbone_bd_ram_mem0_140_0,
         p_wishbone_bd_ram_mem0_140_1, p_wishbone_bd_ram_mem0_140_2,
         p_wishbone_bd_ram_mem0_140_3, p_wishbone_bd_ram_mem0_140_4,
         p_wishbone_bd_ram_mem0_140_5, p_wishbone_bd_ram_mem0_140_6,
         p_wishbone_bd_ram_mem0_140_7, p_wishbone_bd_ram_mem0_141_0,
         p_wishbone_bd_ram_mem0_141_1, p_wishbone_bd_ram_mem0_141_2,
         p_wishbone_bd_ram_mem0_141_3, p_wishbone_bd_ram_mem0_141_4,
         p_wishbone_bd_ram_mem0_141_5, p_wishbone_bd_ram_mem0_141_6,
         p_wishbone_bd_ram_mem0_141_7, p_wishbone_bd_ram_mem0_142_0,
         p_wishbone_bd_ram_mem0_142_1, p_wishbone_bd_ram_mem0_142_2,
         p_wishbone_bd_ram_mem0_142_3, p_wishbone_bd_ram_mem0_142_4,
         p_wishbone_bd_ram_mem0_142_5, p_wishbone_bd_ram_mem0_142_6,
         p_wishbone_bd_ram_mem0_142_7, p_wishbone_bd_ram_mem0_143_0,
         p_wishbone_bd_ram_mem0_143_1, p_wishbone_bd_ram_mem0_143_2,
         p_wishbone_bd_ram_mem0_143_3, p_wishbone_bd_ram_mem0_143_4,
         p_wishbone_bd_ram_mem0_143_5, p_wishbone_bd_ram_mem0_143_6,
         p_wishbone_bd_ram_mem0_143_7, p_wishbone_bd_ram_mem0_144_0,
         p_wishbone_bd_ram_mem0_144_1, p_wishbone_bd_ram_mem0_144_2,
         p_wishbone_bd_ram_mem0_144_3, p_wishbone_bd_ram_mem0_144_4,
         p_wishbone_bd_ram_mem0_144_5, p_wishbone_bd_ram_mem0_144_6,
         p_wishbone_bd_ram_mem0_144_7, p_wishbone_bd_ram_mem0_145_0,
         p_wishbone_bd_ram_mem0_145_1, p_wishbone_bd_ram_mem0_145_2,
         p_wishbone_bd_ram_mem0_145_3, p_wishbone_bd_ram_mem0_145_4,
         p_wishbone_bd_ram_mem0_145_5, p_wishbone_bd_ram_mem0_145_6,
         p_wishbone_bd_ram_mem0_145_7, p_wishbone_bd_ram_mem0_146_0,
         p_wishbone_bd_ram_mem0_146_1, p_wishbone_bd_ram_mem0_146_2,
         p_wishbone_bd_ram_mem0_146_3, p_wishbone_bd_ram_mem0_146_4,
         p_wishbone_bd_ram_mem0_146_5, p_wishbone_bd_ram_mem0_146_6,
         p_wishbone_bd_ram_mem0_146_7, p_wishbone_bd_ram_mem0_147_0,
         p_wishbone_bd_ram_mem0_147_1, p_wishbone_bd_ram_mem0_147_2,
         p_wishbone_bd_ram_mem0_147_3, p_wishbone_bd_ram_mem0_147_4,
         p_wishbone_bd_ram_mem0_147_5, p_wishbone_bd_ram_mem0_147_6,
         p_wishbone_bd_ram_mem0_147_7, p_wishbone_bd_ram_mem0_148_0,
         p_wishbone_bd_ram_mem0_148_1, p_wishbone_bd_ram_mem0_148_2,
         p_wishbone_bd_ram_mem0_148_3, p_wishbone_bd_ram_mem0_148_4,
         p_wishbone_bd_ram_mem0_148_5, p_wishbone_bd_ram_mem0_148_6,
         p_wishbone_bd_ram_mem0_148_7, p_wishbone_bd_ram_mem0_149_0,
         p_wishbone_bd_ram_mem0_149_1, p_wishbone_bd_ram_mem0_149_2,
         p_wishbone_bd_ram_mem0_149_3, p_wishbone_bd_ram_mem0_149_4,
         p_wishbone_bd_ram_mem0_149_5, p_wishbone_bd_ram_mem0_149_6,
         p_wishbone_bd_ram_mem0_149_7, p_wishbone_bd_ram_mem0_150_0,
         p_wishbone_bd_ram_mem0_150_1, p_wishbone_bd_ram_mem0_150_2,
         p_wishbone_bd_ram_mem0_150_3, p_wishbone_bd_ram_mem0_150_4,
         p_wishbone_bd_ram_mem0_150_5, p_wishbone_bd_ram_mem0_150_6,
         p_wishbone_bd_ram_mem0_150_7, p_wishbone_bd_ram_mem0_151_0,
         p_wishbone_bd_ram_mem0_151_1, p_wishbone_bd_ram_mem0_151_2,
         p_wishbone_bd_ram_mem0_151_3, p_wishbone_bd_ram_mem0_151_4,
         p_wishbone_bd_ram_mem0_151_5, p_wishbone_bd_ram_mem0_151_6,
         p_wishbone_bd_ram_mem0_151_7, p_wishbone_bd_ram_mem0_152_0,
         p_wishbone_bd_ram_mem0_152_1, p_wishbone_bd_ram_mem0_152_2,
         p_wishbone_bd_ram_mem0_152_3, p_wishbone_bd_ram_mem0_152_4,
         p_wishbone_bd_ram_mem0_152_5, p_wishbone_bd_ram_mem0_152_6,
         p_wishbone_bd_ram_mem0_152_7, p_wishbone_bd_ram_mem0_153_0,
         p_wishbone_bd_ram_mem0_153_1, p_wishbone_bd_ram_mem0_153_2,
         p_wishbone_bd_ram_mem0_153_3, p_wishbone_bd_ram_mem0_153_4,
         p_wishbone_bd_ram_mem0_153_5, p_wishbone_bd_ram_mem0_153_6,
         p_wishbone_bd_ram_mem0_153_7, p_wishbone_bd_ram_mem0_154_0,
         p_wishbone_bd_ram_mem0_154_1, p_wishbone_bd_ram_mem0_154_2,
         p_wishbone_bd_ram_mem0_154_3, p_wishbone_bd_ram_mem0_154_4,
         p_wishbone_bd_ram_mem0_154_5, p_wishbone_bd_ram_mem0_154_6,
         p_wishbone_bd_ram_mem0_154_7, p_wishbone_bd_ram_mem0_155_0,
         p_wishbone_bd_ram_mem0_155_1, p_wishbone_bd_ram_mem0_155_2,
         p_wishbone_bd_ram_mem0_155_3, p_wishbone_bd_ram_mem0_155_4,
         p_wishbone_bd_ram_mem0_155_5, p_wishbone_bd_ram_mem0_155_6,
         p_wishbone_bd_ram_mem0_155_7, p_wishbone_bd_ram_mem0_156_0,
         p_wishbone_bd_ram_mem0_156_1, p_wishbone_bd_ram_mem0_156_2,
         p_wishbone_bd_ram_mem0_156_3, p_wishbone_bd_ram_mem0_156_4,
         p_wishbone_bd_ram_mem0_156_5, p_wishbone_bd_ram_mem0_156_6,
         p_wishbone_bd_ram_mem0_156_7, p_wishbone_bd_ram_mem0_157_0,
         p_wishbone_bd_ram_mem0_157_1, p_wishbone_bd_ram_mem0_157_2,
         p_wishbone_bd_ram_mem0_157_3, p_wishbone_bd_ram_mem0_157_4,
         p_wishbone_bd_ram_mem0_157_5, p_wishbone_bd_ram_mem0_157_6,
         p_wishbone_bd_ram_mem0_157_7, p_wishbone_bd_ram_mem0_158_0,
         p_wishbone_bd_ram_mem0_158_1, p_wishbone_bd_ram_mem0_158_2,
         p_wishbone_bd_ram_mem0_158_3, p_wishbone_bd_ram_mem0_158_4,
         p_wishbone_bd_ram_mem0_158_5, p_wishbone_bd_ram_mem0_158_6,
         p_wishbone_bd_ram_mem0_158_7, p_wishbone_bd_ram_mem0_159_0,
         p_wishbone_bd_ram_mem0_159_1, p_wishbone_bd_ram_mem0_159_2,
         p_wishbone_bd_ram_mem0_159_3, p_wishbone_bd_ram_mem0_159_4,
         p_wishbone_bd_ram_mem0_159_5, p_wishbone_bd_ram_mem0_159_6,
         p_wishbone_bd_ram_mem0_159_7, p_wishbone_bd_ram_mem0_160_0,
         p_wishbone_bd_ram_mem0_160_1, p_wishbone_bd_ram_mem0_160_2,
         p_wishbone_bd_ram_mem0_160_3, p_wishbone_bd_ram_mem0_160_4,
         p_wishbone_bd_ram_mem0_160_5, p_wishbone_bd_ram_mem0_160_6,
         p_wishbone_bd_ram_mem0_160_7, p_wishbone_bd_ram_mem0_161_0,
         p_wishbone_bd_ram_mem0_161_1, p_wishbone_bd_ram_mem0_161_2,
         p_wishbone_bd_ram_mem0_161_3, p_wishbone_bd_ram_mem0_161_4,
         p_wishbone_bd_ram_mem0_161_5, p_wishbone_bd_ram_mem0_161_6,
         p_wishbone_bd_ram_mem0_161_7, p_wishbone_bd_ram_mem0_162_0,
         p_wishbone_bd_ram_mem0_162_1, p_wishbone_bd_ram_mem0_162_2,
         p_wishbone_bd_ram_mem0_162_3, p_wishbone_bd_ram_mem0_162_4,
         p_wishbone_bd_ram_mem0_162_5, p_wishbone_bd_ram_mem0_162_6,
         p_wishbone_bd_ram_mem0_162_7, p_wishbone_bd_ram_mem0_163_0,
         p_wishbone_bd_ram_mem0_163_1, p_wishbone_bd_ram_mem0_163_2,
         p_wishbone_bd_ram_mem0_163_3, p_wishbone_bd_ram_mem0_163_4,
         p_wishbone_bd_ram_mem0_163_5, p_wishbone_bd_ram_mem0_163_6,
         p_wishbone_bd_ram_mem0_163_7, p_wishbone_bd_ram_mem0_164_0,
         p_wishbone_bd_ram_mem0_164_1, p_wishbone_bd_ram_mem0_164_2,
         p_wishbone_bd_ram_mem0_164_3, p_wishbone_bd_ram_mem0_164_4,
         p_wishbone_bd_ram_mem0_164_5, p_wishbone_bd_ram_mem0_164_6,
         p_wishbone_bd_ram_mem0_164_7, p_wishbone_bd_ram_mem0_165_0,
         p_wishbone_bd_ram_mem0_165_1, p_wishbone_bd_ram_mem0_165_2,
         p_wishbone_bd_ram_mem0_165_3, p_wishbone_bd_ram_mem0_165_4,
         p_wishbone_bd_ram_mem0_165_5, p_wishbone_bd_ram_mem0_165_6,
         p_wishbone_bd_ram_mem0_165_7, p_wishbone_bd_ram_mem0_166_0,
         p_wishbone_bd_ram_mem0_166_1, p_wishbone_bd_ram_mem0_166_2,
         p_wishbone_bd_ram_mem0_166_3, p_wishbone_bd_ram_mem0_166_4,
         p_wishbone_bd_ram_mem0_166_5, p_wishbone_bd_ram_mem0_166_6,
         p_wishbone_bd_ram_mem0_166_7, p_wishbone_bd_ram_mem0_167_0,
         p_wishbone_bd_ram_mem0_167_1, p_wishbone_bd_ram_mem0_167_2,
         p_wishbone_bd_ram_mem0_167_3, p_wishbone_bd_ram_mem0_167_4,
         p_wishbone_bd_ram_mem0_167_5, p_wishbone_bd_ram_mem0_167_6,
         p_wishbone_bd_ram_mem0_167_7, p_wishbone_bd_ram_mem0_168_0,
         p_wishbone_bd_ram_mem0_168_1, p_wishbone_bd_ram_mem0_168_2,
         p_wishbone_bd_ram_mem0_168_3, p_wishbone_bd_ram_mem0_168_4,
         p_wishbone_bd_ram_mem0_168_5, p_wishbone_bd_ram_mem0_168_6,
         p_wishbone_bd_ram_mem0_168_7, p_wishbone_bd_ram_mem0_169_0,
         p_wishbone_bd_ram_mem0_169_1, p_wishbone_bd_ram_mem0_169_2,
         p_wishbone_bd_ram_mem0_169_3, p_wishbone_bd_ram_mem0_169_4,
         p_wishbone_bd_ram_mem0_169_5, p_wishbone_bd_ram_mem0_169_6,
         p_wishbone_bd_ram_mem0_169_7, p_wishbone_bd_ram_mem0_170_0,
         p_wishbone_bd_ram_mem0_170_1, p_wishbone_bd_ram_mem0_170_2,
         p_wishbone_bd_ram_mem0_170_3, p_wishbone_bd_ram_mem0_170_4,
         p_wishbone_bd_ram_mem0_170_5, p_wishbone_bd_ram_mem0_170_6,
         p_wishbone_bd_ram_mem0_170_7, p_wishbone_bd_ram_mem0_171_0,
         p_wishbone_bd_ram_mem0_171_1, p_wishbone_bd_ram_mem0_171_2,
         p_wishbone_bd_ram_mem0_171_3, p_wishbone_bd_ram_mem0_171_4,
         p_wishbone_bd_ram_mem0_171_5, p_wishbone_bd_ram_mem0_171_6,
         p_wishbone_bd_ram_mem0_171_7, p_wishbone_bd_ram_mem0_172_0,
         p_wishbone_bd_ram_mem0_172_1, p_wishbone_bd_ram_mem0_172_2,
         p_wishbone_bd_ram_mem0_172_3, p_wishbone_bd_ram_mem0_172_4,
         p_wishbone_bd_ram_mem0_172_5, p_wishbone_bd_ram_mem0_172_6,
         p_wishbone_bd_ram_mem0_172_7, p_wishbone_bd_ram_mem0_173_0,
         p_wishbone_bd_ram_mem0_173_1, p_wishbone_bd_ram_mem0_173_2,
         p_wishbone_bd_ram_mem0_173_3, p_wishbone_bd_ram_mem0_173_4,
         p_wishbone_bd_ram_mem0_173_5, p_wishbone_bd_ram_mem0_173_6,
         p_wishbone_bd_ram_mem0_173_7, p_wishbone_bd_ram_mem0_174_0,
         p_wishbone_bd_ram_mem0_174_1, p_wishbone_bd_ram_mem0_174_2,
         p_wishbone_bd_ram_mem0_174_3, p_wishbone_bd_ram_mem0_174_4,
         p_wishbone_bd_ram_mem0_174_5, p_wishbone_bd_ram_mem0_174_6,
         p_wishbone_bd_ram_mem0_174_7, p_wishbone_bd_ram_mem0_175_0,
         p_wishbone_bd_ram_mem0_175_1, p_wishbone_bd_ram_mem0_175_2,
         p_wishbone_bd_ram_mem0_175_3, p_wishbone_bd_ram_mem0_175_4,
         p_wishbone_bd_ram_mem0_175_5, p_wishbone_bd_ram_mem0_175_6,
         p_wishbone_bd_ram_mem0_175_7, p_wishbone_bd_ram_mem0_176_0,
         p_wishbone_bd_ram_mem0_176_1, p_wishbone_bd_ram_mem0_176_2,
         p_wishbone_bd_ram_mem0_176_3, p_wishbone_bd_ram_mem0_176_4,
         p_wishbone_bd_ram_mem0_176_5, p_wishbone_bd_ram_mem0_176_6,
         p_wishbone_bd_ram_mem0_176_7, p_wishbone_bd_ram_mem0_177_0,
         p_wishbone_bd_ram_mem0_177_1, p_wishbone_bd_ram_mem0_177_2,
         p_wishbone_bd_ram_mem0_177_3, p_wishbone_bd_ram_mem0_177_4,
         p_wishbone_bd_ram_mem0_177_5, p_wishbone_bd_ram_mem0_177_6,
         p_wishbone_bd_ram_mem0_177_7, p_wishbone_bd_ram_mem0_178_0,
         p_wishbone_bd_ram_mem0_178_1, p_wishbone_bd_ram_mem0_178_2,
         p_wishbone_bd_ram_mem0_178_3, p_wishbone_bd_ram_mem0_178_4,
         p_wishbone_bd_ram_mem0_178_5, p_wishbone_bd_ram_mem0_178_6,
         p_wishbone_bd_ram_mem0_178_7, p_wishbone_bd_ram_mem0_179_0,
         p_wishbone_bd_ram_mem0_179_1, p_wishbone_bd_ram_mem0_179_2,
         p_wishbone_bd_ram_mem0_179_3, p_wishbone_bd_ram_mem0_179_4,
         p_wishbone_bd_ram_mem0_179_5, p_wishbone_bd_ram_mem0_179_6,
         p_wishbone_bd_ram_mem0_179_7, p_wishbone_bd_ram_mem0_180_0,
         p_wishbone_bd_ram_mem0_180_1, p_wishbone_bd_ram_mem0_180_2,
         p_wishbone_bd_ram_mem0_180_3, p_wishbone_bd_ram_mem0_180_4,
         p_wishbone_bd_ram_mem0_180_5, p_wishbone_bd_ram_mem0_180_6,
         p_wishbone_bd_ram_mem0_180_7, p_wishbone_bd_ram_mem0_181_0,
         p_wishbone_bd_ram_mem0_181_1, p_wishbone_bd_ram_mem0_181_2,
         p_wishbone_bd_ram_mem0_181_3, p_wishbone_bd_ram_mem0_181_4,
         p_wishbone_bd_ram_mem0_181_5, p_wishbone_bd_ram_mem0_181_6,
         p_wishbone_bd_ram_mem0_181_7, p_wishbone_bd_ram_mem0_182_0,
         p_wishbone_bd_ram_mem0_182_1, p_wishbone_bd_ram_mem0_182_2,
         p_wishbone_bd_ram_mem0_182_3, p_wishbone_bd_ram_mem0_182_4,
         p_wishbone_bd_ram_mem0_182_5, p_wishbone_bd_ram_mem0_182_6,
         p_wishbone_bd_ram_mem0_182_7, p_wishbone_bd_ram_mem0_183_0,
         p_wishbone_bd_ram_mem0_183_1, p_wishbone_bd_ram_mem0_183_2,
         p_wishbone_bd_ram_mem0_183_3, p_wishbone_bd_ram_mem0_183_4,
         p_wishbone_bd_ram_mem0_183_5, p_wishbone_bd_ram_mem0_183_6,
         p_wishbone_bd_ram_mem0_183_7, p_wishbone_bd_ram_mem0_184_0,
         p_wishbone_bd_ram_mem0_184_1, p_wishbone_bd_ram_mem0_184_2,
         p_wishbone_bd_ram_mem0_184_3, p_wishbone_bd_ram_mem0_184_4,
         p_wishbone_bd_ram_mem0_184_5, p_wishbone_bd_ram_mem0_184_6,
         p_wishbone_bd_ram_mem0_184_7, p_wishbone_bd_ram_mem0_185_0,
         p_wishbone_bd_ram_mem0_185_1, p_wishbone_bd_ram_mem0_185_2,
         p_wishbone_bd_ram_mem0_185_3, p_wishbone_bd_ram_mem0_185_4,
         p_wishbone_bd_ram_mem0_185_5, p_wishbone_bd_ram_mem0_185_6,
         p_wishbone_bd_ram_mem0_185_7, p_wishbone_bd_ram_mem0_186_0,
         p_wishbone_bd_ram_mem0_186_1, p_wishbone_bd_ram_mem0_186_2,
         p_wishbone_bd_ram_mem0_186_3, p_wishbone_bd_ram_mem0_186_4,
         p_wishbone_bd_ram_mem0_186_5, p_wishbone_bd_ram_mem0_186_6,
         p_wishbone_bd_ram_mem0_186_7, p_wishbone_bd_ram_mem0_187_0,
         p_wishbone_bd_ram_mem0_187_1, p_wishbone_bd_ram_mem0_187_2,
         p_wishbone_bd_ram_mem0_187_3, p_wishbone_bd_ram_mem0_187_4,
         p_wishbone_bd_ram_mem0_187_5, p_wishbone_bd_ram_mem0_187_6,
         p_wishbone_bd_ram_mem0_187_7, p_wishbone_bd_ram_mem0_188_0,
         p_wishbone_bd_ram_mem0_188_1, p_wishbone_bd_ram_mem0_188_2,
         p_wishbone_bd_ram_mem0_188_3, p_wishbone_bd_ram_mem0_188_4,
         p_wishbone_bd_ram_mem0_188_5, p_wishbone_bd_ram_mem0_188_6,
         p_wishbone_bd_ram_mem0_188_7, p_wishbone_bd_ram_mem0_189_0,
         p_wishbone_bd_ram_mem0_189_1, p_wishbone_bd_ram_mem0_189_2,
         p_wishbone_bd_ram_mem0_189_3, p_wishbone_bd_ram_mem0_189_4,
         p_wishbone_bd_ram_mem0_189_5, p_wishbone_bd_ram_mem0_189_6,
         p_wishbone_bd_ram_mem0_189_7, p_wishbone_bd_ram_mem0_190_0,
         p_wishbone_bd_ram_mem0_190_1, p_wishbone_bd_ram_mem0_190_2,
         p_wishbone_bd_ram_mem0_190_3, p_wishbone_bd_ram_mem0_190_4,
         p_wishbone_bd_ram_mem0_190_5, p_wishbone_bd_ram_mem0_190_6,
         p_wishbone_bd_ram_mem0_190_7, p_wishbone_bd_ram_mem0_191_0,
         p_wishbone_bd_ram_mem0_191_1, p_wishbone_bd_ram_mem0_191_2,
         p_wishbone_bd_ram_mem0_191_3, p_wishbone_bd_ram_mem0_191_4,
         p_wishbone_bd_ram_mem0_191_5, p_wishbone_bd_ram_mem0_191_6,
         p_wishbone_bd_ram_mem0_191_7, p_wishbone_bd_ram_mem0_192_0,
         p_wishbone_bd_ram_mem0_192_1, p_wishbone_bd_ram_mem0_192_2,
         p_wishbone_bd_ram_mem0_192_3, p_wishbone_bd_ram_mem0_192_4,
         p_wishbone_bd_ram_mem0_192_5, p_wishbone_bd_ram_mem0_192_6,
         p_wishbone_bd_ram_mem0_192_7, p_wishbone_bd_ram_mem0_193_0,
         p_wishbone_bd_ram_mem0_193_1, p_wishbone_bd_ram_mem0_193_2,
         p_wishbone_bd_ram_mem0_193_3, p_wishbone_bd_ram_mem0_193_4,
         p_wishbone_bd_ram_mem0_193_5, p_wishbone_bd_ram_mem0_193_6,
         p_wishbone_bd_ram_mem0_193_7, p_wishbone_bd_ram_mem0_194_0,
         p_wishbone_bd_ram_mem0_194_1, p_wishbone_bd_ram_mem0_194_2,
         p_wishbone_bd_ram_mem0_194_3, p_wishbone_bd_ram_mem0_194_4,
         p_wishbone_bd_ram_mem0_194_5, p_wishbone_bd_ram_mem0_194_6,
         p_wishbone_bd_ram_mem0_194_7, p_wishbone_bd_ram_mem0_195_0,
         p_wishbone_bd_ram_mem0_195_1, p_wishbone_bd_ram_mem0_195_2,
         p_wishbone_bd_ram_mem0_195_3, p_wishbone_bd_ram_mem0_195_4,
         p_wishbone_bd_ram_mem0_195_5, p_wishbone_bd_ram_mem0_195_6,
         p_wishbone_bd_ram_mem0_195_7, p_wishbone_bd_ram_mem0_196_0,
         p_wishbone_bd_ram_mem0_196_1, p_wishbone_bd_ram_mem0_196_2,
         p_wishbone_bd_ram_mem0_196_3, p_wishbone_bd_ram_mem0_196_4,
         p_wishbone_bd_ram_mem0_196_5, p_wishbone_bd_ram_mem0_196_6,
         p_wishbone_bd_ram_mem0_196_7, p_wishbone_bd_ram_mem0_197_0,
         p_wishbone_bd_ram_mem0_197_1, p_wishbone_bd_ram_mem0_197_2,
         p_wishbone_bd_ram_mem0_197_3, p_wishbone_bd_ram_mem0_197_4,
         p_wishbone_bd_ram_mem0_197_5, p_wishbone_bd_ram_mem0_197_6,
         p_wishbone_bd_ram_mem0_197_7, p_wishbone_bd_ram_mem0_198_0,
         p_wishbone_bd_ram_mem0_198_1, p_wishbone_bd_ram_mem0_198_2,
         p_wishbone_bd_ram_mem0_198_3, p_wishbone_bd_ram_mem0_198_4,
         p_wishbone_bd_ram_mem0_198_5, p_wishbone_bd_ram_mem0_198_6,
         p_wishbone_bd_ram_mem0_198_7, p_wishbone_bd_ram_mem0_199_0,
         p_wishbone_bd_ram_mem0_199_1, p_wishbone_bd_ram_mem0_199_2,
         p_wishbone_bd_ram_mem0_199_3, p_wishbone_bd_ram_mem0_199_4,
         p_wishbone_bd_ram_mem0_199_5, p_wishbone_bd_ram_mem0_199_6,
         p_wishbone_bd_ram_mem0_199_7, p_wishbone_bd_ram_mem0_200_0,
         p_wishbone_bd_ram_mem0_200_1, p_wishbone_bd_ram_mem0_200_2,
         p_wishbone_bd_ram_mem0_200_3, p_wishbone_bd_ram_mem0_200_4,
         p_wishbone_bd_ram_mem0_200_5, p_wishbone_bd_ram_mem0_200_6,
         p_wishbone_bd_ram_mem0_200_7, p_wishbone_bd_ram_mem0_201_0,
         p_wishbone_bd_ram_mem0_201_1, p_wishbone_bd_ram_mem0_201_2,
         p_wishbone_bd_ram_mem0_201_3, p_wishbone_bd_ram_mem0_201_4,
         p_wishbone_bd_ram_mem0_201_5, p_wishbone_bd_ram_mem0_201_6,
         p_wishbone_bd_ram_mem0_201_7, p_wishbone_bd_ram_mem0_202_0,
         p_wishbone_bd_ram_mem0_202_1, p_wishbone_bd_ram_mem0_202_2,
         p_wishbone_bd_ram_mem0_202_3, p_wishbone_bd_ram_mem0_202_4,
         p_wishbone_bd_ram_mem0_202_5, p_wishbone_bd_ram_mem0_202_6,
         p_wishbone_bd_ram_mem0_202_7, p_wishbone_bd_ram_mem0_203_0,
         p_wishbone_bd_ram_mem0_203_1, p_wishbone_bd_ram_mem0_203_2,
         p_wishbone_bd_ram_mem0_203_3, p_wishbone_bd_ram_mem0_203_4,
         p_wishbone_bd_ram_mem0_203_5, p_wishbone_bd_ram_mem0_203_6,
         p_wishbone_bd_ram_mem0_203_7, p_wishbone_bd_ram_mem0_204_0,
         p_wishbone_bd_ram_mem0_204_1, p_wishbone_bd_ram_mem0_204_2,
         p_wishbone_bd_ram_mem0_204_3, p_wishbone_bd_ram_mem0_204_4,
         p_wishbone_bd_ram_mem0_204_5, p_wishbone_bd_ram_mem0_204_6,
         p_wishbone_bd_ram_mem0_204_7, p_wishbone_bd_ram_mem0_205_0,
         p_wishbone_bd_ram_mem0_205_1, p_wishbone_bd_ram_mem0_205_2,
         p_wishbone_bd_ram_mem0_205_3, p_wishbone_bd_ram_mem0_205_4,
         p_wishbone_bd_ram_mem0_205_5, p_wishbone_bd_ram_mem0_205_6,
         p_wishbone_bd_ram_mem0_205_7, p_wishbone_bd_ram_mem0_206_0,
         p_wishbone_bd_ram_mem0_206_1, p_wishbone_bd_ram_mem0_206_2,
         p_wishbone_bd_ram_mem0_206_3, p_wishbone_bd_ram_mem0_206_4,
         p_wishbone_bd_ram_mem0_206_5, p_wishbone_bd_ram_mem0_206_6,
         p_wishbone_bd_ram_mem0_206_7, p_wishbone_bd_ram_mem0_207_0,
         p_wishbone_bd_ram_mem0_207_1, p_wishbone_bd_ram_mem0_207_2,
         p_wishbone_bd_ram_mem0_207_3, p_wishbone_bd_ram_mem0_207_4,
         p_wishbone_bd_ram_mem0_207_5, p_wishbone_bd_ram_mem0_207_6,
         p_wishbone_bd_ram_mem0_207_7, p_wishbone_bd_ram_mem0_208_0,
         p_wishbone_bd_ram_mem0_208_1, p_wishbone_bd_ram_mem0_208_2,
         p_wishbone_bd_ram_mem0_208_3, p_wishbone_bd_ram_mem0_208_4,
         p_wishbone_bd_ram_mem0_208_5, p_wishbone_bd_ram_mem0_208_6,
         p_wishbone_bd_ram_mem0_208_7, p_wishbone_bd_ram_mem0_209_0,
         p_wishbone_bd_ram_mem0_209_1, p_wishbone_bd_ram_mem0_209_2,
         p_wishbone_bd_ram_mem0_209_3, p_wishbone_bd_ram_mem0_209_4,
         p_wishbone_bd_ram_mem0_209_5, p_wishbone_bd_ram_mem0_209_6,
         p_wishbone_bd_ram_mem0_209_7, p_wishbone_bd_ram_mem0_210_0,
         p_wishbone_bd_ram_mem0_210_1, p_wishbone_bd_ram_mem0_210_2,
         p_wishbone_bd_ram_mem0_210_3, p_wishbone_bd_ram_mem0_210_4,
         p_wishbone_bd_ram_mem0_210_5, p_wishbone_bd_ram_mem0_210_6,
         p_wishbone_bd_ram_mem0_210_7, p_wishbone_bd_ram_mem0_211_0,
         p_wishbone_bd_ram_mem0_211_1, p_wishbone_bd_ram_mem0_211_2,
         p_wishbone_bd_ram_mem0_211_3, p_wishbone_bd_ram_mem0_211_4,
         p_wishbone_bd_ram_mem0_211_5, p_wishbone_bd_ram_mem0_211_6,
         p_wishbone_bd_ram_mem0_211_7, p_wishbone_bd_ram_mem0_212_0,
         p_wishbone_bd_ram_mem0_212_1, p_wishbone_bd_ram_mem0_212_2,
         p_wishbone_bd_ram_mem0_212_3, p_wishbone_bd_ram_mem0_212_4,
         p_wishbone_bd_ram_mem0_212_5, p_wishbone_bd_ram_mem0_212_6,
         p_wishbone_bd_ram_mem0_212_7, p_wishbone_bd_ram_mem0_213_0,
         p_wishbone_bd_ram_mem0_213_1, p_wishbone_bd_ram_mem0_213_2,
         p_wishbone_bd_ram_mem0_213_3, p_wishbone_bd_ram_mem0_213_4,
         p_wishbone_bd_ram_mem0_213_5, p_wishbone_bd_ram_mem0_213_6,
         p_wishbone_bd_ram_mem0_213_7, p_wishbone_bd_ram_mem0_214_0,
         p_wishbone_bd_ram_mem0_214_1, p_wishbone_bd_ram_mem0_214_2,
         p_wishbone_bd_ram_mem0_214_3, p_wishbone_bd_ram_mem0_214_4,
         p_wishbone_bd_ram_mem0_214_5, p_wishbone_bd_ram_mem0_214_6,
         p_wishbone_bd_ram_mem0_214_7, p_wishbone_bd_ram_mem0_215_0,
         p_wishbone_bd_ram_mem0_215_1, p_wishbone_bd_ram_mem0_215_2,
         p_wishbone_bd_ram_mem0_215_3, p_wishbone_bd_ram_mem0_215_4,
         p_wishbone_bd_ram_mem0_215_5, p_wishbone_bd_ram_mem0_215_6,
         p_wishbone_bd_ram_mem0_215_7, p_wishbone_bd_ram_mem0_216_0,
         p_wishbone_bd_ram_mem0_216_1, p_wishbone_bd_ram_mem0_216_2,
         p_wishbone_bd_ram_mem0_216_3, p_wishbone_bd_ram_mem0_216_4,
         p_wishbone_bd_ram_mem0_216_5, p_wishbone_bd_ram_mem0_216_6,
         p_wishbone_bd_ram_mem0_216_7, p_wishbone_bd_ram_mem0_217_0,
         p_wishbone_bd_ram_mem0_217_1, p_wishbone_bd_ram_mem0_217_2,
         p_wishbone_bd_ram_mem0_217_3, p_wishbone_bd_ram_mem0_217_4,
         p_wishbone_bd_ram_mem0_217_5, p_wishbone_bd_ram_mem0_217_6,
         p_wishbone_bd_ram_mem0_217_7, p_wishbone_bd_ram_mem0_218_0,
         p_wishbone_bd_ram_mem0_218_1, p_wishbone_bd_ram_mem0_218_2,
         p_wishbone_bd_ram_mem0_218_3, p_wishbone_bd_ram_mem0_218_4,
         p_wishbone_bd_ram_mem0_218_5, p_wishbone_bd_ram_mem0_218_6,
         p_wishbone_bd_ram_mem0_218_7, p_wishbone_bd_ram_mem0_219_0,
         p_wishbone_bd_ram_mem0_219_1, p_wishbone_bd_ram_mem0_219_2,
         p_wishbone_bd_ram_mem0_219_3, p_wishbone_bd_ram_mem0_219_4,
         p_wishbone_bd_ram_mem0_219_5, p_wishbone_bd_ram_mem0_219_6,
         p_wishbone_bd_ram_mem0_219_7, p_wishbone_bd_ram_mem0_220_0,
         p_wishbone_bd_ram_mem0_220_1, p_wishbone_bd_ram_mem0_220_2,
         p_wishbone_bd_ram_mem0_220_3, p_wishbone_bd_ram_mem0_220_4,
         p_wishbone_bd_ram_mem0_220_5, p_wishbone_bd_ram_mem0_220_6,
         p_wishbone_bd_ram_mem0_220_7, p_wishbone_bd_ram_mem0_221_0,
         p_wishbone_bd_ram_mem0_221_1, p_wishbone_bd_ram_mem0_221_2,
         p_wishbone_bd_ram_mem0_221_3, p_wishbone_bd_ram_mem0_221_4,
         p_wishbone_bd_ram_mem0_221_5, p_wishbone_bd_ram_mem0_221_6,
         p_wishbone_bd_ram_mem0_221_7, p_wishbone_bd_ram_mem0_222_0,
         p_wishbone_bd_ram_mem0_222_1, p_wishbone_bd_ram_mem0_222_2,
         p_wishbone_bd_ram_mem0_222_3, p_wishbone_bd_ram_mem0_222_4,
         p_wishbone_bd_ram_mem0_222_5, p_wishbone_bd_ram_mem0_222_6,
         p_wishbone_bd_ram_mem0_222_7, p_wishbone_bd_ram_mem0_223_0,
         p_wishbone_bd_ram_mem0_223_1, p_wishbone_bd_ram_mem0_223_2,
         p_wishbone_bd_ram_mem0_223_3, p_wishbone_bd_ram_mem0_223_4,
         p_wishbone_bd_ram_mem0_223_5, p_wishbone_bd_ram_mem0_223_6,
         p_wishbone_bd_ram_mem0_223_7, p_wishbone_bd_ram_mem0_224_0,
         p_wishbone_bd_ram_mem0_224_1, p_wishbone_bd_ram_mem0_224_2,
         p_wishbone_bd_ram_mem0_224_3, p_wishbone_bd_ram_mem0_224_4,
         p_wishbone_bd_ram_mem0_224_5, p_wishbone_bd_ram_mem0_224_6,
         p_wishbone_bd_ram_mem0_224_7, p_wishbone_bd_ram_mem0_225_0,
         p_wishbone_bd_ram_mem0_225_1, p_wishbone_bd_ram_mem0_225_2,
         p_wishbone_bd_ram_mem0_225_3, p_wishbone_bd_ram_mem0_225_4,
         p_wishbone_bd_ram_mem0_225_5, p_wishbone_bd_ram_mem0_225_6,
         p_wishbone_bd_ram_mem0_225_7, p_wishbone_bd_ram_mem0_226_0,
         p_wishbone_bd_ram_mem0_226_1, p_wishbone_bd_ram_mem0_226_2,
         p_wishbone_bd_ram_mem0_226_3, p_wishbone_bd_ram_mem0_226_4,
         p_wishbone_bd_ram_mem0_226_5, p_wishbone_bd_ram_mem0_226_6,
         p_wishbone_bd_ram_mem0_226_7, p_wishbone_bd_ram_mem0_227_0,
         p_wishbone_bd_ram_mem0_227_1, p_wishbone_bd_ram_mem0_227_2,
         p_wishbone_bd_ram_mem0_227_3, p_wishbone_bd_ram_mem0_227_4,
         p_wishbone_bd_ram_mem0_227_5, p_wishbone_bd_ram_mem0_227_6,
         p_wishbone_bd_ram_mem0_227_7, p_wishbone_bd_ram_mem0_228_0,
         p_wishbone_bd_ram_mem0_228_1, p_wishbone_bd_ram_mem0_228_2,
         p_wishbone_bd_ram_mem0_228_3, p_wishbone_bd_ram_mem0_228_4,
         p_wishbone_bd_ram_mem0_228_5, p_wishbone_bd_ram_mem0_228_6,
         p_wishbone_bd_ram_mem0_228_7, p_wishbone_bd_ram_mem0_229_0,
         p_wishbone_bd_ram_mem0_229_1, p_wishbone_bd_ram_mem0_229_2,
         p_wishbone_bd_ram_mem0_229_3, p_wishbone_bd_ram_mem0_229_4,
         p_wishbone_bd_ram_mem0_229_5, p_wishbone_bd_ram_mem0_229_6,
         p_wishbone_bd_ram_mem0_229_7, p_wishbone_bd_ram_mem0_230_0,
         p_wishbone_bd_ram_mem0_230_1, p_wishbone_bd_ram_mem0_230_2,
         p_wishbone_bd_ram_mem0_230_3, p_wishbone_bd_ram_mem0_230_4,
         p_wishbone_bd_ram_mem0_230_5, p_wishbone_bd_ram_mem0_230_6,
         p_wishbone_bd_ram_mem0_230_7, p_wishbone_bd_ram_mem0_231_0,
         p_wishbone_bd_ram_mem0_231_1, p_wishbone_bd_ram_mem0_231_2,
         p_wishbone_bd_ram_mem0_231_3, p_wishbone_bd_ram_mem0_231_4,
         p_wishbone_bd_ram_mem0_231_5, p_wishbone_bd_ram_mem0_231_6,
         p_wishbone_bd_ram_mem0_231_7, p_wishbone_bd_ram_mem0_232_0,
         p_wishbone_bd_ram_mem0_232_1, p_wishbone_bd_ram_mem0_232_2,
         p_wishbone_bd_ram_mem0_232_3, p_wishbone_bd_ram_mem0_232_4,
         p_wishbone_bd_ram_mem0_232_5, p_wishbone_bd_ram_mem0_232_6,
         p_wishbone_bd_ram_mem0_232_7, p_wishbone_bd_ram_mem0_233_0,
         p_wishbone_bd_ram_mem0_233_1, p_wishbone_bd_ram_mem0_233_2,
         p_wishbone_bd_ram_mem0_233_3, p_wishbone_bd_ram_mem0_233_4,
         p_wishbone_bd_ram_mem0_233_5, p_wishbone_bd_ram_mem0_233_6,
         p_wishbone_bd_ram_mem0_233_7, p_wishbone_bd_ram_mem0_234_0,
         p_wishbone_bd_ram_mem0_234_1, p_wishbone_bd_ram_mem0_234_2,
         p_wishbone_bd_ram_mem0_234_3, p_wishbone_bd_ram_mem0_234_4,
         p_wishbone_bd_ram_mem0_234_5, p_wishbone_bd_ram_mem0_234_6,
         p_wishbone_bd_ram_mem0_234_7, p_wishbone_bd_ram_mem0_235_0,
         p_wishbone_bd_ram_mem0_235_1, p_wishbone_bd_ram_mem0_235_2,
         p_wishbone_bd_ram_mem0_235_3, p_wishbone_bd_ram_mem0_235_4,
         p_wishbone_bd_ram_mem0_235_5, p_wishbone_bd_ram_mem0_235_6,
         p_wishbone_bd_ram_mem0_235_7, p_wishbone_bd_ram_mem0_236_0,
         p_wishbone_bd_ram_mem0_236_1, p_wishbone_bd_ram_mem0_236_2,
         p_wishbone_bd_ram_mem0_236_3, p_wishbone_bd_ram_mem0_236_4,
         p_wishbone_bd_ram_mem0_236_5, p_wishbone_bd_ram_mem0_236_6,
         p_wishbone_bd_ram_mem0_236_7, p_wishbone_bd_ram_mem0_237_0,
         p_wishbone_bd_ram_mem0_237_1, p_wishbone_bd_ram_mem0_237_2,
         p_wishbone_bd_ram_mem0_237_3, p_wishbone_bd_ram_mem0_237_4,
         p_wishbone_bd_ram_mem0_237_5, p_wishbone_bd_ram_mem0_237_6,
         p_wishbone_bd_ram_mem0_237_7, p_wishbone_bd_ram_mem0_238_0,
         p_wishbone_bd_ram_mem0_238_1, p_wishbone_bd_ram_mem0_238_2,
         p_wishbone_bd_ram_mem0_238_3, p_wishbone_bd_ram_mem0_238_4,
         p_wishbone_bd_ram_mem0_238_5, p_wishbone_bd_ram_mem0_238_6,
         p_wishbone_bd_ram_mem0_238_7, p_wishbone_bd_ram_mem0_239_0,
         p_wishbone_bd_ram_mem0_239_1, p_wishbone_bd_ram_mem0_239_2,
         p_wishbone_bd_ram_mem0_239_3, p_wishbone_bd_ram_mem0_239_4,
         p_wishbone_bd_ram_mem0_239_5, p_wishbone_bd_ram_mem0_239_6,
         p_wishbone_bd_ram_mem0_239_7, p_wishbone_bd_ram_mem0_240_0,
         p_wishbone_bd_ram_mem0_240_1, p_wishbone_bd_ram_mem0_240_2,
         p_wishbone_bd_ram_mem0_240_3, p_wishbone_bd_ram_mem0_240_4,
         p_wishbone_bd_ram_mem0_240_5, p_wishbone_bd_ram_mem0_240_6,
         p_wishbone_bd_ram_mem0_240_7, p_wishbone_bd_ram_mem0_241_0,
         p_wishbone_bd_ram_mem0_241_1, p_wishbone_bd_ram_mem0_241_2,
         p_wishbone_bd_ram_mem0_241_3, p_wishbone_bd_ram_mem0_241_4,
         p_wishbone_bd_ram_mem0_241_5, p_wishbone_bd_ram_mem0_241_6,
         p_wishbone_bd_ram_mem0_241_7, p_wishbone_bd_ram_mem0_242_0,
         p_wishbone_bd_ram_mem0_242_1, p_wishbone_bd_ram_mem0_242_2,
         p_wishbone_bd_ram_mem0_242_3, p_wishbone_bd_ram_mem0_242_4,
         p_wishbone_bd_ram_mem0_242_5, p_wishbone_bd_ram_mem0_242_6,
         p_wishbone_bd_ram_mem0_242_7, p_wishbone_bd_ram_mem0_243_0,
         p_wishbone_bd_ram_mem0_243_1, p_wishbone_bd_ram_mem0_243_2,
         p_wishbone_bd_ram_mem0_243_3, p_wishbone_bd_ram_mem0_243_4,
         p_wishbone_bd_ram_mem0_243_5, p_wishbone_bd_ram_mem0_243_6,
         p_wishbone_bd_ram_mem0_243_7, p_wishbone_bd_ram_mem0_244_0,
         p_wishbone_bd_ram_mem0_244_1, p_wishbone_bd_ram_mem0_244_2,
         p_wishbone_bd_ram_mem0_244_3, p_wishbone_bd_ram_mem0_244_4,
         p_wishbone_bd_ram_mem0_244_5, p_wishbone_bd_ram_mem0_244_6,
         p_wishbone_bd_ram_mem0_244_7, p_wishbone_bd_ram_mem0_245_0,
         p_wishbone_bd_ram_mem0_245_1, p_wishbone_bd_ram_mem0_245_2,
         p_wishbone_bd_ram_mem0_245_3, p_wishbone_bd_ram_mem0_245_4,
         p_wishbone_bd_ram_mem0_245_5, p_wishbone_bd_ram_mem0_245_6,
         p_wishbone_bd_ram_mem0_245_7, p_wishbone_bd_ram_mem0_246_0,
         p_wishbone_bd_ram_mem0_246_1, p_wishbone_bd_ram_mem0_246_2,
         p_wishbone_bd_ram_mem0_246_3, p_wishbone_bd_ram_mem0_246_4,
         p_wishbone_bd_ram_mem0_246_5, p_wishbone_bd_ram_mem0_246_6,
         p_wishbone_bd_ram_mem0_246_7, p_wishbone_bd_ram_mem0_247_0,
         p_wishbone_bd_ram_mem0_247_1, p_wishbone_bd_ram_mem0_247_2,
         p_wishbone_bd_ram_mem0_247_3, p_wishbone_bd_ram_mem0_247_4,
         p_wishbone_bd_ram_mem0_247_5, p_wishbone_bd_ram_mem0_247_6,
         p_wishbone_bd_ram_mem0_247_7, p_wishbone_bd_ram_mem0_248_0,
         p_wishbone_bd_ram_mem0_248_1, p_wishbone_bd_ram_mem0_248_2,
         p_wishbone_bd_ram_mem0_248_3, p_wishbone_bd_ram_mem0_248_4,
         p_wishbone_bd_ram_mem0_248_5, p_wishbone_bd_ram_mem0_248_6,
         p_wishbone_bd_ram_mem0_248_7, p_wishbone_bd_ram_mem0_249_0,
         p_wishbone_bd_ram_mem0_249_1, p_wishbone_bd_ram_mem0_249_2,
         p_wishbone_bd_ram_mem0_249_3, p_wishbone_bd_ram_mem0_249_4,
         p_wishbone_bd_ram_mem0_249_5, p_wishbone_bd_ram_mem0_249_6,
         p_wishbone_bd_ram_mem0_249_7, p_wishbone_bd_ram_mem0_250_0,
         p_wishbone_bd_ram_mem0_250_1, p_wishbone_bd_ram_mem0_250_2,
         p_wishbone_bd_ram_mem0_250_3, p_wishbone_bd_ram_mem0_250_4,
         p_wishbone_bd_ram_mem0_250_5, p_wishbone_bd_ram_mem0_250_6,
         p_wishbone_bd_ram_mem0_250_7, p_wishbone_bd_ram_mem0_251_0,
         p_wishbone_bd_ram_mem0_251_1, p_wishbone_bd_ram_mem0_251_2,
         p_wishbone_bd_ram_mem0_251_3, p_wishbone_bd_ram_mem0_251_4,
         p_wishbone_bd_ram_mem0_251_5, p_wishbone_bd_ram_mem0_251_6,
         p_wishbone_bd_ram_mem0_251_7, p_wishbone_bd_ram_mem0_252_0,
         p_wishbone_bd_ram_mem0_252_1, p_wishbone_bd_ram_mem0_252_2,
         p_wishbone_bd_ram_mem0_252_3, p_wishbone_bd_ram_mem0_252_4,
         p_wishbone_bd_ram_mem0_252_5, p_wishbone_bd_ram_mem0_252_6,
         p_wishbone_bd_ram_mem0_252_7, p_wishbone_bd_ram_mem0_253_0,
         p_wishbone_bd_ram_mem0_253_1, p_wishbone_bd_ram_mem0_253_2,
         p_wishbone_bd_ram_mem0_253_3, p_wishbone_bd_ram_mem0_253_4,
         p_wishbone_bd_ram_mem0_253_5, p_wishbone_bd_ram_mem0_253_6,
         p_wishbone_bd_ram_mem0_253_7, p_wishbone_bd_ram_mem0_254_0,
         p_wishbone_bd_ram_mem0_254_1, p_wishbone_bd_ram_mem0_254_2,
         p_wishbone_bd_ram_mem0_254_3, p_wishbone_bd_ram_mem0_254_4,
         p_wishbone_bd_ram_mem0_254_5, p_wishbone_bd_ram_mem0_254_6,
         p_wishbone_bd_ram_mem0_254_7, p_wishbone_bd_ram_mem0_255_0,
         p_wishbone_bd_ram_mem0_255_1, p_wishbone_bd_ram_mem0_255_2,
         p_wishbone_bd_ram_mem0_255_3, p_wishbone_bd_ram_mem0_255_4,
         p_wishbone_bd_ram_mem0_255_5, p_wishbone_bd_ram_mem0_255_6,
         p_wishbone_bd_ram_mem0_255_7, p_wishbone_bd_ram_N102,
         p_wishbone_bd_ram_N103, p_wishbone_bd_ram_N104,
         p_wishbone_bd_ram_N105, p_wishbone_bd_ram_N106,
         p_wishbone_bd_ram_N107, p_wishbone_bd_ram_N108,
         p_wishbone_bd_ram_N109, p_wishbone_TxData_wb_0,
         p_wishbone_TxData_wb_1, p_wishbone_TxData_wb_2,
         p_wishbone_TxData_wb_3, p_wishbone_TxData_wb_4,
         p_wishbone_TxData_wb_5, p_wishbone_TxData_wb_6,
         p_wishbone_TxData_wb_7, p_wishbone_TxData_wb_8,
         p_wishbone_TxData_wb_9, p_wishbone_TxData_wb_10,
         p_wishbone_TxData_wb_11, p_wishbone_TxData_wb_12,
         p_wishbone_TxData_wb_13, p_wishbone_TxData_wb_14,
         p_wishbone_TxData_wb_15, p_wishbone_TxData_wb_16,
         p_wishbone_TxData_wb_17, p_wishbone_TxData_wb_18,
         p_wishbone_TxData_wb_19, p_wishbone_TxData_wb_20,
         p_wishbone_TxData_wb_21, p_wishbone_TxData_wb_22,
         p_wishbone_TxData_wb_23, p_wishbone_TxData_wb_24,
         p_wishbone_TxData_wb_25, p_wishbone_TxData_wb_26,
         p_wishbone_TxData_wb_27, p_wishbone_TxData_wb_28,
         p_wishbone_TxData_wb_29, p_wishbone_TxData_wb_30,
         p_wishbone_TxData_wb_31, p_wishbone_tx_fifo_fifo_15_0,
         p_wishbone_tx_fifo_fifo_15_1, p_wishbone_tx_fifo_fifo_15_2,
         p_wishbone_tx_fifo_fifo_15_3, p_wishbone_tx_fifo_fifo_15_4,
         p_wishbone_tx_fifo_fifo_15_5, p_wishbone_tx_fifo_fifo_15_6,
         p_wishbone_tx_fifo_fifo_15_7, p_wishbone_tx_fifo_fifo_15_8,
         p_wishbone_tx_fifo_fifo_15_9, p_wishbone_tx_fifo_fifo_15_10,
         p_wishbone_tx_fifo_fifo_15_11, p_wishbone_tx_fifo_fifo_15_12,
         p_wishbone_tx_fifo_fifo_15_13, p_wishbone_tx_fifo_fifo_15_14,
         p_wishbone_tx_fifo_fifo_15_15, p_wishbone_tx_fifo_fifo_15_16,
         p_wishbone_tx_fifo_fifo_15_17, p_wishbone_tx_fifo_fifo_15_18,
         p_wishbone_tx_fifo_fifo_15_19, p_wishbone_tx_fifo_fifo_15_20,
         p_wishbone_tx_fifo_fifo_15_21, p_wishbone_tx_fifo_fifo_15_22,
         p_wishbone_tx_fifo_fifo_15_23, p_wishbone_tx_fifo_fifo_15_24,
         p_wishbone_tx_fifo_fifo_15_25, p_wishbone_tx_fifo_fifo_15_26,
         p_wishbone_tx_fifo_fifo_15_27, p_wishbone_tx_fifo_fifo_15_28,
         p_wishbone_tx_fifo_fifo_15_29, p_wishbone_tx_fifo_fifo_15_30,
         p_wishbone_tx_fifo_fifo_15_31, p_wishbone_tx_fifo_fifo_14_0,
         p_wishbone_tx_fifo_fifo_14_1, p_wishbone_tx_fifo_fifo_14_2,
         p_wishbone_tx_fifo_fifo_14_3, p_wishbone_tx_fifo_fifo_14_4,
         p_wishbone_tx_fifo_fifo_14_5, p_wishbone_tx_fifo_fifo_14_6,
         p_wishbone_tx_fifo_fifo_14_7, p_wishbone_tx_fifo_fifo_14_8,
         p_wishbone_tx_fifo_fifo_14_9, p_wishbone_tx_fifo_fifo_14_10,
         p_wishbone_tx_fifo_fifo_14_11, p_wishbone_tx_fifo_fifo_14_12,
         p_wishbone_tx_fifo_fifo_14_13, p_wishbone_tx_fifo_fifo_14_14,
         p_wishbone_tx_fifo_fifo_14_15, p_wishbone_tx_fifo_fifo_14_16,
         p_wishbone_tx_fifo_fifo_14_17, p_wishbone_tx_fifo_fifo_14_18,
         p_wishbone_tx_fifo_fifo_14_19, p_wishbone_tx_fifo_fifo_14_20,
         p_wishbone_tx_fifo_fifo_14_21, p_wishbone_tx_fifo_fifo_14_22,
         p_wishbone_tx_fifo_fifo_14_23, p_wishbone_tx_fifo_fifo_14_24,
         p_wishbone_tx_fifo_fifo_14_25, p_wishbone_tx_fifo_fifo_14_26,
         p_wishbone_tx_fifo_fifo_14_27, p_wishbone_tx_fifo_fifo_14_28,
         p_wishbone_tx_fifo_fifo_14_29, p_wishbone_tx_fifo_fifo_14_30,
         p_wishbone_tx_fifo_fifo_14_31, p_wishbone_tx_fifo_fifo_13_0,
         p_wishbone_tx_fifo_fifo_13_1, p_wishbone_tx_fifo_fifo_13_2,
         p_wishbone_tx_fifo_fifo_13_3, p_wishbone_tx_fifo_fifo_13_4,
         p_wishbone_tx_fifo_fifo_13_5, p_wishbone_tx_fifo_fifo_13_6,
         p_wishbone_tx_fifo_fifo_13_7, p_wishbone_tx_fifo_fifo_13_8,
         p_wishbone_tx_fifo_fifo_13_9, p_wishbone_tx_fifo_fifo_13_10,
         p_wishbone_tx_fifo_fifo_13_11, p_wishbone_tx_fifo_fifo_13_12,
         p_wishbone_tx_fifo_fifo_13_13, p_wishbone_tx_fifo_fifo_13_14,
         p_wishbone_tx_fifo_fifo_13_15, p_wishbone_tx_fifo_fifo_13_16,
         p_wishbone_tx_fifo_fifo_13_17, p_wishbone_tx_fifo_fifo_13_18,
         p_wishbone_tx_fifo_fifo_13_19, p_wishbone_tx_fifo_fifo_13_20,
         p_wishbone_tx_fifo_fifo_13_21, p_wishbone_tx_fifo_fifo_13_22,
         p_wishbone_tx_fifo_fifo_13_23, p_wishbone_tx_fifo_fifo_13_24,
         p_wishbone_tx_fifo_fifo_13_25, p_wishbone_tx_fifo_fifo_13_26,
         p_wishbone_tx_fifo_fifo_13_27, p_wishbone_tx_fifo_fifo_13_28,
         p_wishbone_tx_fifo_fifo_13_29, p_wishbone_tx_fifo_fifo_13_30,
         p_wishbone_tx_fifo_fifo_13_31, p_wishbone_tx_fifo_fifo_12_0,
         p_wishbone_tx_fifo_fifo_12_1, p_wishbone_tx_fifo_fifo_12_2,
         p_wishbone_tx_fifo_fifo_12_3, p_wishbone_tx_fifo_fifo_12_4,
         p_wishbone_tx_fifo_fifo_12_5, p_wishbone_tx_fifo_fifo_12_6,
         p_wishbone_tx_fifo_fifo_12_7, p_wishbone_tx_fifo_fifo_12_8,
         p_wishbone_tx_fifo_fifo_12_9, p_wishbone_tx_fifo_fifo_12_10,
         p_wishbone_tx_fifo_fifo_12_11, p_wishbone_tx_fifo_fifo_12_12,
         p_wishbone_tx_fifo_fifo_12_13, p_wishbone_tx_fifo_fifo_12_14,
         p_wishbone_tx_fifo_fifo_12_15, p_wishbone_tx_fifo_fifo_12_16,
         p_wishbone_tx_fifo_fifo_12_17, p_wishbone_tx_fifo_fifo_12_18,
         p_wishbone_tx_fifo_fifo_12_19, p_wishbone_tx_fifo_fifo_12_20,
         p_wishbone_tx_fifo_fifo_12_21, p_wishbone_tx_fifo_fifo_12_22,
         p_wishbone_tx_fifo_fifo_12_23, p_wishbone_tx_fifo_fifo_12_24,
         p_wishbone_tx_fifo_fifo_12_25, p_wishbone_tx_fifo_fifo_12_26,
         p_wishbone_tx_fifo_fifo_12_27, p_wishbone_tx_fifo_fifo_12_28,
         p_wishbone_tx_fifo_fifo_12_29, p_wishbone_tx_fifo_fifo_12_30,
         p_wishbone_tx_fifo_fifo_12_31, p_wishbone_tx_fifo_fifo_11_0,
         p_wishbone_tx_fifo_fifo_11_1, p_wishbone_tx_fifo_fifo_11_2,
         p_wishbone_tx_fifo_fifo_11_3, p_wishbone_tx_fifo_fifo_11_4,
         p_wishbone_tx_fifo_fifo_11_5, p_wishbone_tx_fifo_fifo_11_6,
         p_wishbone_tx_fifo_fifo_11_7, p_wishbone_tx_fifo_fifo_11_8,
         p_wishbone_tx_fifo_fifo_11_9, p_wishbone_tx_fifo_fifo_11_10,
         p_wishbone_tx_fifo_fifo_11_11, p_wishbone_tx_fifo_fifo_11_12,
         p_wishbone_tx_fifo_fifo_11_13, p_wishbone_tx_fifo_fifo_11_14,
         p_wishbone_tx_fifo_fifo_11_15, p_wishbone_tx_fifo_fifo_11_16,
         p_wishbone_tx_fifo_fifo_11_17, p_wishbone_tx_fifo_fifo_11_18,
         p_wishbone_tx_fifo_fifo_11_19, p_wishbone_tx_fifo_fifo_11_20,
         p_wishbone_tx_fifo_fifo_11_21, p_wishbone_tx_fifo_fifo_11_22,
         p_wishbone_tx_fifo_fifo_11_23, p_wishbone_tx_fifo_fifo_11_24,
         p_wishbone_tx_fifo_fifo_11_25, p_wishbone_tx_fifo_fifo_11_26,
         p_wishbone_tx_fifo_fifo_11_27, p_wishbone_tx_fifo_fifo_11_28,
         p_wishbone_tx_fifo_fifo_11_29, p_wishbone_tx_fifo_fifo_11_30,
         p_wishbone_tx_fifo_fifo_11_31, p_wishbone_tx_fifo_fifo_10_0,
         p_wishbone_tx_fifo_fifo_10_1, p_wishbone_tx_fifo_fifo_10_2,
         p_wishbone_tx_fifo_fifo_10_3, p_wishbone_tx_fifo_fifo_10_4,
         p_wishbone_tx_fifo_fifo_10_5, p_wishbone_tx_fifo_fifo_10_6,
         p_wishbone_tx_fifo_fifo_10_7, p_wishbone_tx_fifo_fifo_10_8,
         p_wishbone_tx_fifo_fifo_10_9, p_wishbone_tx_fifo_fifo_10_10,
         p_wishbone_tx_fifo_fifo_10_11, p_wishbone_tx_fifo_fifo_10_12,
         p_wishbone_tx_fifo_fifo_10_13, p_wishbone_tx_fifo_fifo_10_14,
         p_wishbone_tx_fifo_fifo_10_15, p_wishbone_tx_fifo_fifo_10_16,
         p_wishbone_tx_fifo_fifo_10_17, p_wishbone_tx_fifo_fifo_10_18,
         p_wishbone_tx_fifo_fifo_10_19, p_wishbone_tx_fifo_fifo_10_20,
         p_wishbone_tx_fifo_fifo_10_21, p_wishbone_tx_fifo_fifo_10_22,
         p_wishbone_tx_fifo_fifo_10_23, p_wishbone_tx_fifo_fifo_10_24,
         p_wishbone_tx_fifo_fifo_10_25, p_wishbone_tx_fifo_fifo_10_26,
         p_wishbone_tx_fifo_fifo_10_27, p_wishbone_tx_fifo_fifo_10_28,
         p_wishbone_tx_fifo_fifo_10_29, p_wishbone_tx_fifo_fifo_10_30,
         p_wishbone_tx_fifo_fifo_10_31, p_wishbone_tx_fifo_fifo_9_0,
         p_wishbone_tx_fifo_fifo_9_1, p_wishbone_tx_fifo_fifo_9_2,
         p_wishbone_tx_fifo_fifo_9_3, p_wishbone_tx_fifo_fifo_9_4,
         p_wishbone_tx_fifo_fifo_9_5, p_wishbone_tx_fifo_fifo_9_6,
         p_wishbone_tx_fifo_fifo_9_7, p_wishbone_tx_fifo_fifo_9_8,
         p_wishbone_tx_fifo_fifo_9_9, p_wishbone_tx_fifo_fifo_9_10,
         p_wishbone_tx_fifo_fifo_9_11, p_wishbone_tx_fifo_fifo_9_12,
         p_wishbone_tx_fifo_fifo_9_13, p_wishbone_tx_fifo_fifo_9_14,
         p_wishbone_tx_fifo_fifo_9_15, p_wishbone_tx_fifo_fifo_9_16,
         p_wishbone_tx_fifo_fifo_9_17, p_wishbone_tx_fifo_fifo_9_18,
         p_wishbone_tx_fifo_fifo_9_19, p_wishbone_tx_fifo_fifo_9_20,
         p_wishbone_tx_fifo_fifo_9_21, p_wishbone_tx_fifo_fifo_9_22,
         p_wishbone_tx_fifo_fifo_9_23, p_wishbone_tx_fifo_fifo_9_24,
         p_wishbone_tx_fifo_fifo_9_25, p_wishbone_tx_fifo_fifo_9_26,
         p_wishbone_tx_fifo_fifo_9_27, p_wishbone_tx_fifo_fifo_9_28,
         p_wishbone_tx_fifo_fifo_9_29, p_wishbone_tx_fifo_fifo_9_30,
         p_wishbone_tx_fifo_fifo_9_31, p_wishbone_tx_fifo_fifo_8_0,
         p_wishbone_tx_fifo_fifo_8_1, p_wishbone_tx_fifo_fifo_8_2,
         p_wishbone_tx_fifo_fifo_8_3, p_wishbone_tx_fifo_fifo_8_4,
         p_wishbone_tx_fifo_fifo_8_5, p_wishbone_tx_fifo_fifo_8_6,
         p_wishbone_tx_fifo_fifo_8_7, p_wishbone_tx_fifo_fifo_8_8,
         p_wishbone_tx_fifo_fifo_8_9, p_wishbone_tx_fifo_fifo_8_10,
         p_wishbone_tx_fifo_fifo_8_11, p_wishbone_tx_fifo_fifo_8_12,
         p_wishbone_tx_fifo_fifo_8_13, p_wishbone_tx_fifo_fifo_8_14,
         p_wishbone_tx_fifo_fifo_8_15, p_wishbone_tx_fifo_fifo_8_16,
         p_wishbone_tx_fifo_fifo_8_17, p_wishbone_tx_fifo_fifo_8_18,
         p_wishbone_tx_fifo_fifo_8_19, p_wishbone_tx_fifo_fifo_8_20,
         p_wishbone_tx_fifo_fifo_8_21, p_wishbone_tx_fifo_fifo_8_22,
         p_wishbone_tx_fifo_fifo_8_23, p_wishbone_tx_fifo_fifo_8_24,
         p_wishbone_tx_fifo_fifo_8_25, p_wishbone_tx_fifo_fifo_8_26,
         p_wishbone_tx_fifo_fifo_8_27, p_wishbone_tx_fifo_fifo_8_28,
         p_wishbone_tx_fifo_fifo_8_29, p_wishbone_tx_fifo_fifo_8_30,
         p_wishbone_tx_fifo_fifo_8_31, p_wishbone_tx_fifo_fifo_7_0,
         p_wishbone_tx_fifo_fifo_7_1, p_wishbone_tx_fifo_fifo_7_2,
         p_wishbone_tx_fifo_fifo_7_3, p_wishbone_tx_fifo_fifo_7_4,
         p_wishbone_tx_fifo_fifo_7_5, p_wishbone_tx_fifo_fifo_7_6,
         p_wishbone_tx_fifo_fifo_7_7, p_wishbone_tx_fifo_fifo_7_8,
         p_wishbone_tx_fifo_fifo_7_9, p_wishbone_tx_fifo_fifo_7_10,
         p_wishbone_tx_fifo_fifo_7_11, p_wishbone_tx_fifo_fifo_7_12,
         p_wishbone_tx_fifo_fifo_7_13, p_wishbone_tx_fifo_fifo_7_14,
         p_wishbone_tx_fifo_fifo_7_15, p_wishbone_tx_fifo_fifo_7_16,
         p_wishbone_tx_fifo_fifo_7_17, p_wishbone_tx_fifo_fifo_7_18,
         p_wishbone_tx_fifo_fifo_7_19, p_wishbone_tx_fifo_fifo_7_20,
         p_wishbone_tx_fifo_fifo_7_21, p_wishbone_tx_fifo_fifo_7_22,
         p_wishbone_tx_fifo_fifo_7_23, p_wishbone_tx_fifo_fifo_7_24,
         p_wishbone_tx_fifo_fifo_7_25, p_wishbone_tx_fifo_fifo_7_26,
         p_wishbone_tx_fifo_fifo_7_27, p_wishbone_tx_fifo_fifo_7_28,
         p_wishbone_tx_fifo_fifo_7_29, p_wishbone_tx_fifo_fifo_7_30,
         p_wishbone_tx_fifo_fifo_7_31, p_wishbone_tx_fifo_fifo_6_0,
         p_wishbone_tx_fifo_fifo_6_1, p_wishbone_tx_fifo_fifo_6_2,
         p_wishbone_tx_fifo_fifo_6_3, p_wishbone_tx_fifo_fifo_6_4,
         p_wishbone_tx_fifo_fifo_6_5, p_wishbone_tx_fifo_fifo_6_6,
         p_wishbone_tx_fifo_fifo_6_7, p_wishbone_tx_fifo_fifo_6_8,
         p_wishbone_tx_fifo_fifo_6_9, p_wishbone_tx_fifo_fifo_6_10,
         p_wishbone_tx_fifo_fifo_6_11, p_wishbone_tx_fifo_fifo_6_12,
         p_wishbone_tx_fifo_fifo_6_13, p_wishbone_tx_fifo_fifo_6_14,
         p_wishbone_tx_fifo_fifo_6_15, p_wishbone_tx_fifo_fifo_6_16,
         p_wishbone_tx_fifo_fifo_6_17, p_wishbone_tx_fifo_fifo_6_18,
         p_wishbone_tx_fifo_fifo_6_19, p_wishbone_tx_fifo_fifo_6_20,
         p_wishbone_tx_fifo_fifo_6_21, p_wishbone_tx_fifo_fifo_6_22,
         p_wishbone_tx_fifo_fifo_6_23, p_wishbone_tx_fifo_fifo_6_24,
         p_wishbone_tx_fifo_fifo_6_25, p_wishbone_tx_fifo_fifo_6_26,
         p_wishbone_tx_fifo_fifo_6_27, p_wishbone_tx_fifo_fifo_6_28,
         p_wishbone_tx_fifo_fifo_6_29, p_wishbone_tx_fifo_fifo_6_30,
         p_wishbone_tx_fifo_fifo_6_31, p_wishbone_tx_fifo_fifo_5_0,
         p_wishbone_tx_fifo_fifo_5_1, p_wishbone_tx_fifo_fifo_5_2,
         p_wishbone_tx_fifo_fifo_5_3, p_wishbone_tx_fifo_fifo_5_4,
         p_wishbone_tx_fifo_fifo_5_5, p_wishbone_tx_fifo_fifo_5_6,
         p_wishbone_tx_fifo_fifo_5_7, p_wishbone_tx_fifo_fifo_5_8,
         p_wishbone_tx_fifo_fifo_5_9, p_wishbone_tx_fifo_fifo_5_10,
         p_wishbone_tx_fifo_fifo_5_11, p_wishbone_tx_fifo_fifo_5_12,
         p_wishbone_tx_fifo_fifo_5_13, p_wishbone_tx_fifo_fifo_5_14,
         p_wishbone_tx_fifo_fifo_5_15, p_wishbone_tx_fifo_fifo_5_16,
         p_wishbone_tx_fifo_fifo_5_17, p_wishbone_tx_fifo_fifo_5_18,
         p_wishbone_tx_fifo_fifo_5_19, p_wishbone_tx_fifo_fifo_5_20,
         p_wishbone_tx_fifo_fifo_5_21, p_wishbone_tx_fifo_fifo_5_22,
         p_wishbone_tx_fifo_fifo_5_23, p_wishbone_tx_fifo_fifo_5_24,
         p_wishbone_tx_fifo_fifo_5_25, p_wishbone_tx_fifo_fifo_5_26,
         p_wishbone_tx_fifo_fifo_5_27, p_wishbone_tx_fifo_fifo_5_28,
         p_wishbone_tx_fifo_fifo_5_29, p_wishbone_tx_fifo_fifo_5_30,
         p_wishbone_tx_fifo_fifo_5_31, p_wishbone_tx_fifo_fifo_4_0,
         p_wishbone_tx_fifo_fifo_4_1, p_wishbone_tx_fifo_fifo_4_2,
         p_wishbone_tx_fifo_fifo_4_3, p_wishbone_tx_fifo_fifo_4_4,
         p_wishbone_tx_fifo_fifo_4_5, p_wishbone_tx_fifo_fifo_4_6,
         p_wishbone_tx_fifo_fifo_4_7, p_wishbone_tx_fifo_fifo_4_8,
         p_wishbone_tx_fifo_fifo_4_9, p_wishbone_tx_fifo_fifo_4_10,
         p_wishbone_tx_fifo_fifo_4_11, p_wishbone_tx_fifo_fifo_4_12,
         p_wishbone_tx_fifo_fifo_4_13, p_wishbone_tx_fifo_fifo_4_14,
         p_wishbone_tx_fifo_fifo_4_15, p_wishbone_tx_fifo_fifo_4_16,
         p_wishbone_tx_fifo_fifo_4_17, p_wishbone_tx_fifo_fifo_4_18,
         p_wishbone_tx_fifo_fifo_4_19, p_wishbone_tx_fifo_fifo_4_20,
         p_wishbone_tx_fifo_fifo_4_21, p_wishbone_tx_fifo_fifo_4_22,
         p_wishbone_tx_fifo_fifo_4_23, p_wishbone_tx_fifo_fifo_4_24,
         p_wishbone_tx_fifo_fifo_4_25, p_wishbone_tx_fifo_fifo_4_26,
         p_wishbone_tx_fifo_fifo_4_27, p_wishbone_tx_fifo_fifo_4_28,
         p_wishbone_tx_fifo_fifo_4_29, p_wishbone_tx_fifo_fifo_4_30,
         p_wishbone_tx_fifo_fifo_4_31, p_wishbone_tx_fifo_fifo_3_0,
         p_wishbone_tx_fifo_fifo_3_1, p_wishbone_tx_fifo_fifo_3_2,
         p_wishbone_tx_fifo_fifo_3_3, p_wishbone_tx_fifo_fifo_3_4,
         p_wishbone_tx_fifo_fifo_3_5, p_wishbone_tx_fifo_fifo_3_6,
         p_wishbone_tx_fifo_fifo_3_7, p_wishbone_tx_fifo_fifo_3_8,
         p_wishbone_tx_fifo_fifo_3_9, p_wishbone_tx_fifo_fifo_3_10,
         p_wishbone_tx_fifo_fifo_3_11, p_wishbone_tx_fifo_fifo_3_12,
         p_wishbone_tx_fifo_fifo_3_13, p_wishbone_tx_fifo_fifo_3_14,
         p_wishbone_tx_fifo_fifo_3_15, p_wishbone_tx_fifo_fifo_3_16,
         p_wishbone_tx_fifo_fifo_3_17, p_wishbone_tx_fifo_fifo_3_18,
         p_wishbone_tx_fifo_fifo_3_19, p_wishbone_tx_fifo_fifo_3_20,
         p_wishbone_tx_fifo_fifo_3_21, p_wishbone_tx_fifo_fifo_3_22,
         p_wishbone_tx_fifo_fifo_3_23, p_wishbone_tx_fifo_fifo_3_24,
         p_wishbone_tx_fifo_fifo_3_25, p_wishbone_tx_fifo_fifo_3_26,
         p_wishbone_tx_fifo_fifo_3_27, p_wishbone_tx_fifo_fifo_3_28,
         p_wishbone_tx_fifo_fifo_3_29, p_wishbone_tx_fifo_fifo_3_30,
         p_wishbone_tx_fifo_fifo_3_31, p_wishbone_tx_fifo_fifo_2_0,
         p_wishbone_tx_fifo_fifo_2_1, p_wishbone_tx_fifo_fifo_2_2,
         p_wishbone_tx_fifo_fifo_2_3, p_wishbone_tx_fifo_fifo_2_4,
         p_wishbone_tx_fifo_fifo_2_5, p_wishbone_tx_fifo_fifo_2_6,
         p_wishbone_tx_fifo_fifo_2_7, p_wishbone_tx_fifo_fifo_2_8,
         p_wishbone_tx_fifo_fifo_2_9, p_wishbone_tx_fifo_fifo_2_10,
         p_wishbone_tx_fifo_fifo_2_11, p_wishbone_tx_fifo_fifo_2_12,
         p_wishbone_tx_fifo_fifo_2_13, p_wishbone_tx_fifo_fifo_2_14,
         p_wishbone_tx_fifo_fifo_2_15, p_wishbone_tx_fifo_fifo_2_16,
         p_wishbone_tx_fifo_fifo_2_17, p_wishbone_tx_fifo_fifo_2_18,
         p_wishbone_tx_fifo_fifo_2_19, p_wishbone_tx_fifo_fifo_2_20,
         p_wishbone_tx_fifo_fifo_2_21, p_wishbone_tx_fifo_fifo_2_22,
         p_wishbone_tx_fifo_fifo_2_23, p_wishbone_tx_fifo_fifo_2_24,
         p_wishbone_tx_fifo_fifo_2_25, p_wishbone_tx_fifo_fifo_2_26,
         p_wishbone_tx_fifo_fifo_2_27, p_wishbone_tx_fifo_fifo_2_28,
         p_wishbone_tx_fifo_fifo_2_29, p_wishbone_tx_fifo_fifo_2_30,
         p_wishbone_tx_fifo_fifo_2_31, p_wishbone_tx_fifo_fifo_1_0,
         p_wishbone_tx_fifo_fifo_1_1, p_wishbone_tx_fifo_fifo_1_2,
         p_wishbone_tx_fifo_fifo_1_3, p_wishbone_tx_fifo_fifo_1_4,
         p_wishbone_tx_fifo_fifo_1_5, p_wishbone_tx_fifo_fifo_1_6,
         p_wishbone_tx_fifo_fifo_1_7, p_wishbone_tx_fifo_fifo_1_8,
         p_wishbone_tx_fifo_fifo_1_9, p_wishbone_tx_fifo_fifo_1_10,
         p_wishbone_tx_fifo_fifo_1_11, p_wishbone_tx_fifo_fifo_1_12,
         p_wishbone_tx_fifo_fifo_1_13, p_wishbone_tx_fifo_fifo_1_14,
         p_wishbone_tx_fifo_fifo_1_15, p_wishbone_tx_fifo_fifo_1_16,
         p_wishbone_tx_fifo_fifo_1_17, p_wishbone_tx_fifo_fifo_1_18,
         p_wishbone_tx_fifo_fifo_1_19, p_wishbone_tx_fifo_fifo_1_20,
         p_wishbone_tx_fifo_fifo_1_21, p_wishbone_tx_fifo_fifo_1_22,
         p_wishbone_tx_fifo_fifo_1_23, p_wishbone_tx_fifo_fifo_1_24,
         p_wishbone_tx_fifo_fifo_1_25, p_wishbone_tx_fifo_fifo_1_26,
         p_wishbone_tx_fifo_fifo_1_27, p_wishbone_tx_fifo_fifo_1_28,
         p_wishbone_tx_fifo_fifo_1_29, p_wishbone_tx_fifo_fifo_1_30,
         p_wishbone_tx_fifo_fifo_1_31, p_wishbone_tx_fifo_fifo_0_0,
         p_wishbone_tx_fifo_fifo_0_1, p_wishbone_tx_fifo_fifo_0_2,
         p_wishbone_tx_fifo_fifo_0_3, p_wishbone_tx_fifo_fifo_0_4,
         p_wishbone_tx_fifo_fifo_0_5, p_wishbone_tx_fifo_fifo_0_6,
         p_wishbone_tx_fifo_fifo_0_7, p_wishbone_tx_fifo_fifo_0_8,
         p_wishbone_tx_fifo_fifo_0_9, p_wishbone_tx_fifo_fifo_0_10,
         p_wishbone_tx_fifo_fifo_0_11, p_wishbone_tx_fifo_fifo_0_12,
         p_wishbone_tx_fifo_fifo_0_13, p_wishbone_tx_fifo_fifo_0_14,
         p_wishbone_tx_fifo_fifo_0_15, p_wishbone_tx_fifo_fifo_0_16,
         p_wishbone_tx_fifo_fifo_0_17, p_wishbone_tx_fifo_fifo_0_18,
         p_wishbone_tx_fifo_fifo_0_19, p_wishbone_tx_fifo_fifo_0_20,
         p_wishbone_tx_fifo_fifo_0_21, p_wishbone_tx_fifo_fifo_0_22,
         p_wishbone_tx_fifo_fifo_0_23, p_wishbone_tx_fifo_fifo_0_24,
         p_wishbone_tx_fifo_fifo_0_25, p_wishbone_tx_fifo_fifo_0_26,
         p_wishbone_tx_fifo_fifo_0_27, p_wishbone_tx_fifo_fifo_0_28,
         p_wishbone_tx_fifo_fifo_0_29, p_wishbone_tx_fifo_fifo_0_30,
         p_wishbone_tx_fifo_fifo_0_31, p_wishbone_tx_fifo_write_pointer_3,
         p_wishbone_tx_fifo_write_pointer_2,
         p_wishbone_tx_fifo_write_pointer_1,
         p_wishbone_tx_fifo_write_pointer_0, p_wishbone_tx_fifo_N17,
         p_wishbone_tx_fifo_N16, p_wishbone_tx_fifo_N15,
         p_wishbone_tx_fifo_N14, p_wishbone_txfifo_cnt_4,
         p_wishbone_txfifo_cnt_3, p_wishbone_txfifo_cnt_2,
         p_wishbone_txfifo_cnt_1, p_wishbone_txfifo_cnt_0, r_TxPauseTV_8,
         r_TxPauseTV_9, r_TxPauseTV_10, r_TxPauseTV_11, r_TxPauseTV_12,
         r_TxPauseTV_13, r_TxPauseTV_14, r_TxPauseTV_15, r_TxPauseTV_0,
         r_TxPauseTV_1, r_TxPauseTV_2, r_TxPauseTV_3, r_TxPauseTV_4,
         r_TxPauseTV_5, r_TxPauseTV_6, r_TxPauseTV_7, r_HASH1_24, r_HASH1_25,
         r_HASH1_26, r_HASH1_27, r_HASH1_28, r_HASH1_29, r_HASH1_30,
         r_HASH1_31, r_HASH1_16, r_HASH1_17, r_HASH1_18, r_HASH1_19,
         r_HASH1_20, r_HASH1_21, r_HASH1_22, r_HASH1_23, r_HASH1_8, r_HASH1_9,
         r_HASH1_10, r_HASH1_11, r_HASH1_12, r_HASH1_13, r_HASH1_14,
         r_HASH1_15, r_HASH1_0, r_HASH1_1, r_HASH1_2, r_HASH1_3, r_HASH1_4,
         r_HASH1_5, r_HASH1_6, r_HASH1_7, r_HASH0_24, r_HASH0_25, r_HASH0_26,
         r_HASH0_27, r_HASH0_28, r_HASH0_29, r_HASH0_30, r_HASH0_31,
         r_HASH0_16, r_HASH0_17, r_HASH0_18, r_HASH0_19, r_HASH0_20,
         r_HASH0_21, r_HASH0_22, r_HASH0_23, r_HASH0_8, r_HASH0_9, r_HASH0_10,
         r_HASH0_11, r_HASH0_12, r_HASH0_13, r_HASH0_14, r_HASH0_15, r_HASH0_0,
         r_HASH0_1, r_HASH0_2, r_HASH0_3, r_HASH0_4, r_HASH0_5, r_HASH0_6,
         r_HASH0_7, r_MAC_40, r_MAC_41, r_MAC_42, r_MAC_43, r_MAC_44, r_MAC_45,
         r_MAC_46, r_MAC_47, r_MAC_32, r_MAC_33, r_MAC_34, r_MAC_35, r_MAC_36,
         r_MAC_37, r_MAC_38, r_MAC_39, r_MAC_24, r_MAC_25, r_MAC_26, r_MAC_27,
         r_MAC_28, r_MAC_29, r_MAC_30, r_MAC_31, r_MAC_16, r_MAC_17, r_MAC_18,
         r_MAC_19, r_MAC_20, r_MAC_21, r_MAC_22, r_MAC_23, r_MAC_8, r_MAC_9,
         r_MAC_10, r_MAC_11, r_MAC_12, r_MAC_13, r_MAC_14, r_MAC_15, r_MAC_0,
         r_MAC_1, r_MAC_2, r_MAC_3, r_MAC_4, r_MAC_5, r_MAC_6, r_MAC_7,
         r_CtrlData_8, r_CtrlData_9, r_CtrlData_10, r_CtrlData_11,
         r_CtrlData_12, r_CtrlData_13, r_CtrlData_14, r_CtrlData_15,
         r_CtrlData_0, r_CtrlData_1, r_CtrlData_2, r_CtrlData_3, r_CtrlData_4,
         r_CtrlData_5, r_CtrlData_6, r_CtrlData_7, r_MinFL_8, r_MinFL_9,
         r_MinFL_10, r_MinFL_11, r_MinFL_12, r_MinFL_13, r_MinFL_14,
         r_MinFL_15, r_MaxFL_0, r_MaxFL_1, r_MaxFL_2, r_MaxFL_3, r_MaxFL_4,
         r_MaxFL_5, r_MaxFL_6, r_MaxFL_7, r_TxPauseRq, r_MiiNoPre, r_IPGR2_0,
         r_IPGR2_1, r_IPGR2_2, r_IPGR2_3, r_IPGR2_4, r_IPGR2_5, r_IPGR2_6,
         r_TxBDNum_0, r_TxBDNum_1, r_TxBDNum_2, r_TxBDNum_3, r_TxBDNum_4,
         r_TxBDNum_5, r_TxBDNum_6, r_TxBDNum_7, r_RGAD_0, r_RGAD_1, r_RGAD_2,
         r_RGAD_3, r_RGAD_4, p_rxethmac1_crcrx_Crc_22,
         p_rxethmac1_crcrx_Crc_18, p_rxethmac1_crcrx_Crc_14,
         p_rxethmac1_crcrx_Crc_10, p_rxethmac1_crcrx_Crc_6,
         p_rxethmac1_crcrx_Crc_2, p_rxethmac1_crcrx_Crc_5,
         p_rxethmac1_crcrx_Crc_23, p_rxethmac1_crcrx_Crc_19,
         p_rxethmac1_crcrx_Crc_15, p_rxethmac1_crcrx_Crc_11,
         p_rxethmac1_crcrx_Crc_7, p_rxethmac1_crcrx_Crc_3, p_rxethmac1_Crc_31,
         p_rxethmac1_Crc_27, p_rxethmac1_crcrx_Crc_1, p_rxethmac1_Crc_29,
         p_rxethmac1_crcrx_Crc_25, p_rxethmac1_crcrx_Crc_21,
         p_rxethmac1_crcrx_Crc_17, p_rxethmac1_crcrx_Crc_13,
         p_rxethmac1_crcrx_Crc_9, p_rxethmac1_Crc_30, p_rxethmac1_Crc_26,
         p_rxethmac1_Crc_28, p_rxethmac1_crcrx_Crc_24,
         p_rxethmac1_crcrx_Crc_20, p_rxethmac1_crcrx_Crc_16,
         p_rxethmac1_crcrx_Crc_12, p_rxethmac1_crcrx_Crc_8,
         p_rxethmac1_crcrx_Crc_4, p_rxethmac1_crcrx_Crc_0,
         p_wishbone_rx_fifo_fifo_15_0, p_wishbone_rx_fifo_fifo_15_1,
         p_wishbone_rx_fifo_fifo_15_2, p_wishbone_rx_fifo_fifo_15_3,
         p_wishbone_rx_fifo_fifo_15_4, p_wishbone_rx_fifo_fifo_15_5,
         p_wishbone_rx_fifo_fifo_15_6, p_wishbone_rx_fifo_fifo_15_7,
         p_wishbone_rx_fifo_fifo_15_8, p_wishbone_rx_fifo_fifo_15_9,
         p_wishbone_rx_fifo_fifo_15_10, p_wishbone_rx_fifo_fifo_15_11,
         p_wishbone_rx_fifo_fifo_15_12, p_wishbone_rx_fifo_fifo_15_13,
         p_wishbone_rx_fifo_fifo_15_14, p_wishbone_rx_fifo_fifo_15_15,
         p_wishbone_rx_fifo_fifo_15_16, p_wishbone_rx_fifo_fifo_15_17,
         p_wishbone_rx_fifo_fifo_15_18, p_wishbone_rx_fifo_fifo_15_19,
         p_wishbone_rx_fifo_fifo_15_20, p_wishbone_rx_fifo_fifo_15_21,
         p_wishbone_rx_fifo_fifo_15_22, p_wishbone_rx_fifo_fifo_15_23,
         p_wishbone_rx_fifo_fifo_15_24, p_wishbone_rx_fifo_fifo_15_25,
         p_wishbone_rx_fifo_fifo_15_26, p_wishbone_rx_fifo_fifo_15_27,
         p_wishbone_rx_fifo_fifo_15_28, p_wishbone_rx_fifo_fifo_15_29,
         p_wishbone_rx_fifo_fifo_15_30, p_wishbone_rx_fifo_fifo_15_31,
         p_wishbone_rx_fifo_fifo_14_0, p_wishbone_rx_fifo_fifo_14_1,
         p_wishbone_rx_fifo_fifo_14_2, p_wishbone_rx_fifo_fifo_14_3,
         p_wishbone_rx_fifo_fifo_14_4, p_wishbone_rx_fifo_fifo_14_5,
         p_wishbone_rx_fifo_fifo_14_6, p_wishbone_rx_fifo_fifo_14_7,
         p_wishbone_rx_fifo_fifo_14_8, p_wishbone_rx_fifo_fifo_14_9,
         p_wishbone_rx_fifo_fifo_14_10, p_wishbone_rx_fifo_fifo_14_11,
         p_wishbone_rx_fifo_fifo_14_12, p_wishbone_rx_fifo_fifo_14_13,
         p_wishbone_rx_fifo_fifo_14_14, p_wishbone_rx_fifo_fifo_14_15,
         p_wishbone_rx_fifo_fifo_14_16, p_wishbone_rx_fifo_fifo_14_17,
         p_wishbone_rx_fifo_fifo_14_18, p_wishbone_rx_fifo_fifo_14_19,
         p_wishbone_rx_fifo_fifo_14_20, p_wishbone_rx_fifo_fifo_14_21,
         p_wishbone_rx_fifo_fifo_14_22, p_wishbone_rx_fifo_fifo_14_23,
         p_wishbone_rx_fifo_fifo_14_24, p_wishbone_rx_fifo_fifo_14_25,
         p_wishbone_rx_fifo_fifo_14_26, p_wishbone_rx_fifo_fifo_14_27,
         p_wishbone_rx_fifo_fifo_14_28, p_wishbone_rx_fifo_fifo_14_29,
         p_wishbone_rx_fifo_fifo_14_30, p_wishbone_rx_fifo_fifo_14_31,
         p_wishbone_rx_fifo_fifo_13_0, p_wishbone_rx_fifo_fifo_13_1,
         p_wishbone_rx_fifo_fifo_13_2, p_wishbone_rx_fifo_fifo_13_3,
         p_wishbone_rx_fifo_fifo_13_4, p_wishbone_rx_fifo_fifo_13_5,
         p_wishbone_rx_fifo_fifo_13_6, p_wishbone_rx_fifo_fifo_13_7,
         p_wishbone_rx_fifo_fifo_13_8, p_wishbone_rx_fifo_fifo_13_9,
         p_wishbone_rx_fifo_fifo_13_10, p_wishbone_rx_fifo_fifo_13_11,
         p_wishbone_rx_fifo_fifo_13_12, p_wishbone_rx_fifo_fifo_13_13,
         p_wishbone_rx_fifo_fifo_13_14, p_wishbone_rx_fifo_fifo_13_15,
         p_wishbone_rx_fifo_fifo_13_16, p_wishbone_rx_fifo_fifo_13_17,
         p_wishbone_rx_fifo_fifo_13_18, p_wishbone_rx_fifo_fifo_13_19,
         p_wishbone_rx_fifo_fifo_13_20, p_wishbone_rx_fifo_fifo_13_21,
         p_wishbone_rx_fifo_fifo_13_22, p_wishbone_rx_fifo_fifo_13_23,
         p_wishbone_rx_fifo_fifo_13_24, p_wishbone_rx_fifo_fifo_13_25,
         p_wishbone_rx_fifo_fifo_13_26, p_wishbone_rx_fifo_fifo_13_27,
         p_wishbone_rx_fifo_fifo_13_28, p_wishbone_rx_fifo_fifo_13_29,
         p_wishbone_rx_fifo_fifo_13_30, p_wishbone_rx_fifo_fifo_13_31,
         p_wishbone_rx_fifo_fifo_12_0, p_wishbone_rx_fifo_fifo_12_1,
         p_wishbone_rx_fifo_fifo_12_2, p_wishbone_rx_fifo_fifo_12_3,
         p_wishbone_rx_fifo_fifo_12_4, p_wishbone_rx_fifo_fifo_12_5,
         p_wishbone_rx_fifo_fifo_12_6, p_wishbone_rx_fifo_fifo_12_7,
         p_wishbone_rx_fifo_fifo_12_8, p_wishbone_rx_fifo_fifo_12_9,
         p_wishbone_rx_fifo_fifo_12_10, p_wishbone_rx_fifo_fifo_12_11,
         p_wishbone_rx_fifo_fifo_12_12, p_wishbone_rx_fifo_fifo_12_13,
         p_wishbone_rx_fifo_fifo_12_14, p_wishbone_rx_fifo_fifo_12_15,
         p_wishbone_rx_fifo_fifo_12_16, p_wishbone_rx_fifo_fifo_12_17,
         p_wishbone_rx_fifo_fifo_12_18, p_wishbone_rx_fifo_fifo_12_19,
         p_wishbone_rx_fifo_fifo_12_20, p_wishbone_rx_fifo_fifo_12_21,
         p_wishbone_rx_fifo_fifo_12_22, p_wishbone_rx_fifo_fifo_12_23,
         p_wishbone_rx_fifo_fifo_12_24, p_wishbone_rx_fifo_fifo_12_25,
         p_wishbone_rx_fifo_fifo_12_26, p_wishbone_rx_fifo_fifo_12_27,
         p_wishbone_rx_fifo_fifo_12_28, p_wishbone_rx_fifo_fifo_12_29,
         p_wishbone_rx_fifo_fifo_12_30, p_wishbone_rx_fifo_fifo_12_31,
         p_wishbone_rx_fifo_fifo_11_0, p_wishbone_rx_fifo_fifo_11_1,
         p_wishbone_rx_fifo_fifo_11_2, p_wishbone_rx_fifo_fifo_11_3,
         p_wishbone_rx_fifo_fifo_11_4, p_wishbone_rx_fifo_fifo_11_5,
         p_wishbone_rx_fifo_fifo_11_6, p_wishbone_rx_fifo_fifo_11_7,
         p_wishbone_rx_fifo_fifo_11_8, p_wishbone_rx_fifo_fifo_11_9,
         p_wishbone_rx_fifo_fifo_11_10, p_wishbone_rx_fifo_fifo_11_11,
         p_wishbone_rx_fifo_fifo_11_12, p_wishbone_rx_fifo_fifo_11_13,
         p_wishbone_rx_fifo_fifo_11_14, p_wishbone_rx_fifo_fifo_11_15,
         p_wishbone_rx_fifo_fifo_11_16, p_wishbone_rx_fifo_fifo_11_17,
         p_wishbone_rx_fifo_fifo_11_18, p_wishbone_rx_fifo_fifo_11_19,
         p_wishbone_rx_fifo_fifo_11_20, p_wishbone_rx_fifo_fifo_11_21,
         p_wishbone_rx_fifo_fifo_11_22, p_wishbone_rx_fifo_fifo_11_23,
         p_wishbone_rx_fifo_fifo_11_24, p_wishbone_rx_fifo_fifo_11_25,
         p_wishbone_rx_fifo_fifo_11_26, p_wishbone_rx_fifo_fifo_11_27,
         p_wishbone_rx_fifo_fifo_11_28, p_wishbone_rx_fifo_fifo_11_29,
         p_wishbone_rx_fifo_fifo_11_30, p_wishbone_rx_fifo_fifo_11_31,
         p_wishbone_rx_fifo_fifo_10_0, p_wishbone_rx_fifo_fifo_10_1,
         p_wishbone_rx_fifo_fifo_10_2, p_wishbone_rx_fifo_fifo_10_3,
         p_wishbone_rx_fifo_fifo_10_4, p_wishbone_rx_fifo_fifo_10_5,
         p_wishbone_rx_fifo_fifo_10_6, p_wishbone_rx_fifo_fifo_10_7,
         p_wishbone_rx_fifo_fifo_10_8, p_wishbone_rx_fifo_fifo_10_9,
         p_wishbone_rx_fifo_fifo_10_10, p_wishbone_rx_fifo_fifo_10_11,
         p_wishbone_rx_fifo_fifo_10_12, p_wishbone_rx_fifo_fifo_10_13,
         p_wishbone_rx_fifo_fifo_10_14, p_wishbone_rx_fifo_fifo_10_15,
         p_wishbone_rx_fifo_fifo_10_16, p_wishbone_rx_fifo_fifo_10_17,
         p_wishbone_rx_fifo_fifo_10_18, p_wishbone_rx_fifo_fifo_10_19,
         p_wishbone_rx_fifo_fifo_10_20, p_wishbone_rx_fifo_fifo_10_21,
         p_wishbone_rx_fifo_fifo_10_22, p_wishbone_rx_fifo_fifo_10_23,
         p_wishbone_rx_fifo_fifo_10_24, p_wishbone_rx_fifo_fifo_10_25,
         p_wishbone_rx_fifo_fifo_10_26, p_wishbone_rx_fifo_fifo_10_27,
         p_wishbone_rx_fifo_fifo_10_28, p_wishbone_rx_fifo_fifo_10_29,
         p_wishbone_rx_fifo_fifo_10_30, p_wishbone_rx_fifo_fifo_10_31,
         p_wishbone_rx_fifo_fifo_9_0, p_wishbone_rx_fifo_fifo_9_1,
         p_wishbone_rx_fifo_fifo_9_2, p_wishbone_rx_fifo_fifo_9_3,
         p_wishbone_rx_fifo_fifo_9_4, p_wishbone_rx_fifo_fifo_9_5,
         p_wishbone_rx_fifo_fifo_9_6, p_wishbone_rx_fifo_fifo_9_7,
         p_wishbone_rx_fifo_fifo_9_8, p_wishbone_rx_fifo_fifo_9_9,
         p_wishbone_rx_fifo_fifo_9_10, p_wishbone_rx_fifo_fifo_9_11,
         p_wishbone_rx_fifo_fifo_9_12, p_wishbone_rx_fifo_fifo_9_13,
         p_wishbone_rx_fifo_fifo_9_14, p_wishbone_rx_fifo_fifo_9_15,
         p_wishbone_rx_fifo_fifo_9_16, p_wishbone_rx_fifo_fifo_9_17,
         p_wishbone_rx_fifo_fifo_9_18, p_wishbone_rx_fifo_fifo_9_19,
         p_wishbone_rx_fifo_fifo_9_20, p_wishbone_rx_fifo_fifo_9_21,
         p_wishbone_rx_fifo_fifo_9_22, p_wishbone_rx_fifo_fifo_9_23,
         p_wishbone_rx_fifo_fifo_9_24, p_wishbone_rx_fifo_fifo_9_25,
         p_wishbone_rx_fifo_fifo_9_26, p_wishbone_rx_fifo_fifo_9_27,
         p_wishbone_rx_fifo_fifo_9_28, p_wishbone_rx_fifo_fifo_9_29,
         p_wishbone_rx_fifo_fifo_9_30, p_wishbone_rx_fifo_fifo_9_31,
         p_wishbone_rx_fifo_fifo_8_0, p_wishbone_rx_fifo_fifo_8_1,
         p_wishbone_rx_fifo_fifo_8_2, p_wishbone_rx_fifo_fifo_8_3,
         p_wishbone_rx_fifo_fifo_8_4, p_wishbone_rx_fifo_fifo_8_5,
         p_wishbone_rx_fifo_fifo_8_6, p_wishbone_rx_fifo_fifo_8_7,
         p_wishbone_rx_fifo_fifo_8_8, p_wishbone_rx_fifo_fifo_8_9,
         p_wishbone_rx_fifo_fifo_8_10, p_wishbone_rx_fifo_fifo_8_11,
         p_wishbone_rx_fifo_fifo_8_12, p_wishbone_rx_fifo_fifo_8_13,
         p_wishbone_rx_fifo_fifo_8_14, p_wishbone_rx_fifo_fifo_8_15,
         p_wishbone_rx_fifo_fifo_8_16, p_wishbone_rx_fifo_fifo_8_17,
         p_wishbone_rx_fifo_fifo_8_18, p_wishbone_rx_fifo_fifo_8_19,
         p_wishbone_rx_fifo_fifo_8_20, p_wishbone_rx_fifo_fifo_8_21,
         p_wishbone_rx_fifo_fifo_8_22, p_wishbone_rx_fifo_fifo_8_23,
         p_wishbone_rx_fifo_fifo_8_24, p_wishbone_rx_fifo_fifo_8_25,
         p_wishbone_rx_fifo_fifo_8_26, p_wishbone_rx_fifo_fifo_8_27,
         p_wishbone_rx_fifo_fifo_8_28, p_wishbone_rx_fifo_fifo_8_29,
         p_wishbone_rx_fifo_fifo_8_30, p_wishbone_rx_fifo_fifo_8_31,
         p_wishbone_rx_fifo_fifo_7_0, p_wishbone_rx_fifo_fifo_7_1,
         p_wishbone_rx_fifo_fifo_7_2, p_wishbone_rx_fifo_fifo_7_3,
         p_wishbone_rx_fifo_fifo_7_4, p_wishbone_rx_fifo_fifo_7_5,
         p_wishbone_rx_fifo_fifo_7_6, p_wishbone_rx_fifo_fifo_7_7,
         p_wishbone_rx_fifo_fifo_7_8, p_wishbone_rx_fifo_fifo_7_9,
         p_wishbone_rx_fifo_fifo_7_10, p_wishbone_rx_fifo_fifo_7_11,
         p_wishbone_rx_fifo_fifo_7_12, p_wishbone_rx_fifo_fifo_7_13,
         p_wishbone_rx_fifo_fifo_7_14, p_wishbone_rx_fifo_fifo_7_15,
         p_wishbone_rx_fifo_fifo_7_16, p_wishbone_rx_fifo_fifo_7_17,
         p_wishbone_rx_fifo_fifo_7_18, p_wishbone_rx_fifo_fifo_7_19,
         p_wishbone_rx_fifo_fifo_7_20, p_wishbone_rx_fifo_fifo_7_21,
         p_wishbone_rx_fifo_fifo_7_22, p_wishbone_rx_fifo_fifo_7_23,
         p_wishbone_rx_fifo_fifo_7_24, p_wishbone_rx_fifo_fifo_7_25,
         p_wishbone_rx_fifo_fifo_7_26, p_wishbone_rx_fifo_fifo_7_27,
         p_wishbone_rx_fifo_fifo_7_28, p_wishbone_rx_fifo_fifo_7_29,
         p_wishbone_rx_fifo_fifo_7_30, p_wishbone_rx_fifo_fifo_7_31,
         p_wishbone_rx_fifo_fifo_6_0, p_wishbone_rx_fifo_fifo_6_1,
         p_wishbone_rx_fifo_fifo_6_2, p_wishbone_rx_fifo_fifo_6_3,
         p_wishbone_rx_fifo_fifo_6_4, p_wishbone_rx_fifo_fifo_6_5,
         p_wishbone_rx_fifo_fifo_6_6, p_wishbone_rx_fifo_fifo_6_7,
         p_wishbone_rx_fifo_fifo_6_8, p_wishbone_rx_fifo_fifo_6_9,
         p_wishbone_rx_fifo_fifo_6_10, p_wishbone_rx_fifo_fifo_6_11,
         p_wishbone_rx_fifo_fifo_6_12, p_wishbone_rx_fifo_fifo_6_13,
         p_wishbone_rx_fifo_fifo_6_14, p_wishbone_rx_fifo_fifo_6_15,
         p_wishbone_rx_fifo_fifo_6_16, p_wishbone_rx_fifo_fifo_6_17,
         p_wishbone_rx_fifo_fifo_6_18, p_wishbone_rx_fifo_fifo_6_19,
         p_wishbone_rx_fifo_fifo_6_20, p_wishbone_rx_fifo_fifo_6_21,
         p_wishbone_rx_fifo_fifo_6_22, p_wishbone_rx_fifo_fifo_6_23,
         p_wishbone_rx_fifo_fifo_6_24, p_wishbone_rx_fifo_fifo_6_25,
         p_wishbone_rx_fifo_fifo_6_26, p_wishbone_rx_fifo_fifo_6_27,
         p_wishbone_rx_fifo_fifo_6_28, p_wishbone_rx_fifo_fifo_6_29,
         p_wishbone_rx_fifo_fifo_6_30, p_wishbone_rx_fifo_fifo_6_31,
         p_wishbone_rx_fifo_fifo_5_0, p_wishbone_rx_fifo_fifo_5_1,
         p_wishbone_rx_fifo_fifo_5_2, p_wishbone_rx_fifo_fifo_5_3,
         p_wishbone_rx_fifo_fifo_5_4, p_wishbone_rx_fifo_fifo_5_5,
         p_wishbone_rx_fifo_fifo_5_6, p_wishbone_rx_fifo_fifo_5_7,
         p_wishbone_rx_fifo_fifo_5_8, p_wishbone_rx_fifo_fifo_5_9,
         p_wishbone_rx_fifo_fifo_5_10, p_wishbone_rx_fifo_fifo_5_11,
         p_wishbone_rx_fifo_fifo_5_12, p_wishbone_rx_fifo_fifo_5_13,
         p_wishbone_rx_fifo_fifo_5_14, p_wishbone_rx_fifo_fifo_5_15,
         p_wishbone_rx_fifo_fifo_5_16, p_wishbone_rx_fifo_fifo_5_17,
         p_wishbone_rx_fifo_fifo_5_18, p_wishbone_rx_fifo_fifo_5_19,
         p_wishbone_rx_fifo_fifo_5_20, p_wishbone_rx_fifo_fifo_5_21,
         p_wishbone_rx_fifo_fifo_5_22, p_wishbone_rx_fifo_fifo_5_23,
         p_wishbone_rx_fifo_fifo_5_24, p_wishbone_rx_fifo_fifo_5_25,
         p_wishbone_rx_fifo_fifo_5_26, p_wishbone_rx_fifo_fifo_5_27,
         p_wishbone_rx_fifo_fifo_5_28, p_wishbone_rx_fifo_fifo_5_29,
         p_wishbone_rx_fifo_fifo_5_30, p_wishbone_rx_fifo_fifo_5_31,
         p_wishbone_rx_fifo_fifo_4_0, p_wishbone_rx_fifo_fifo_4_1,
         p_wishbone_rx_fifo_fifo_4_2, p_wishbone_rx_fifo_fifo_4_3,
         p_wishbone_rx_fifo_fifo_4_4, p_wishbone_rx_fifo_fifo_4_5,
         p_wishbone_rx_fifo_fifo_4_6, p_wishbone_rx_fifo_fifo_4_7,
         p_wishbone_rx_fifo_fifo_4_8, p_wishbone_rx_fifo_fifo_4_9,
         p_wishbone_rx_fifo_fifo_4_10, p_wishbone_rx_fifo_fifo_4_11,
         p_wishbone_rx_fifo_fifo_4_12, p_wishbone_rx_fifo_fifo_4_13,
         p_wishbone_rx_fifo_fifo_4_14, p_wishbone_rx_fifo_fifo_4_15,
         p_wishbone_rx_fifo_fifo_4_16, p_wishbone_rx_fifo_fifo_4_17,
         p_wishbone_rx_fifo_fifo_4_18, p_wishbone_rx_fifo_fifo_4_19,
         p_wishbone_rx_fifo_fifo_4_20, p_wishbone_rx_fifo_fifo_4_21,
         p_wishbone_rx_fifo_fifo_4_22, p_wishbone_rx_fifo_fifo_4_23,
         p_wishbone_rx_fifo_fifo_4_24, p_wishbone_rx_fifo_fifo_4_25,
         p_wishbone_rx_fifo_fifo_4_26, p_wishbone_rx_fifo_fifo_4_27,
         p_wishbone_rx_fifo_fifo_4_28, p_wishbone_rx_fifo_fifo_4_29,
         p_wishbone_rx_fifo_fifo_4_30, p_wishbone_rx_fifo_fifo_4_31,
         p_wishbone_rx_fifo_fifo_3_0, p_wishbone_rx_fifo_fifo_3_1,
         p_wishbone_rx_fifo_fifo_3_2, p_wishbone_rx_fifo_fifo_3_3,
         p_wishbone_rx_fifo_fifo_3_4, p_wishbone_rx_fifo_fifo_3_5,
         p_wishbone_rx_fifo_fifo_3_6, p_wishbone_rx_fifo_fifo_3_7,
         p_wishbone_rx_fifo_fifo_3_8, p_wishbone_rx_fifo_fifo_3_9,
         p_wishbone_rx_fifo_fifo_3_10, p_wishbone_rx_fifo_fifo_3_11,
         p_wishbone_rx_fifo_fifo_3_12, p_wishbone_rx_fifo_fifo_3_13,
         p_wishbone_rx_fifo_fifo_3_14, p_wishbone_rx_fifo_fifo_3_15,
         p_wishbone_rx_fifo_fifo_3_16, p_wishbone_rx_fifo_fifo_3_17,
         p_wishbone_rx_fifo_fifo_3_18, p_wishbone_rx_fifo_fifo_3_19,
         p_wishbone_rx_fifo_fifo_3_20, p_wishbone_rx_fifo_fifo_3_21,
         p_wishbone_rx_fifo_fifo_3_22, p_wishbone_rx_fifo_fifo_3_23,
         p_wishbone_rx_fifo_fifo_3_24, p_wishbone_rx_fifo_fifo_3_25,
         p_wishbone_rx_fifo_fifo_3_26, p_wishbone_rx_fifo_fifo_3_27,
         p_wishbone_rx_fifo_fifo_3_28, p_wishbone_rx_fifo_fifo_3_29,
         p_wishbone_rx_fifo_fifo_3_30, p_wishbone_rx_fifo_fifo_3_31,
         p_wishbone_rx_fifo_fifo_2_0, p_wishbone_rx_fifo_fifo_2_1,
         p_wishbone_rx_fifo_fifo_2_2, p_wishbone_rx_fifo_fifo_2_3,
         p_wishbone_rx_fifo_fifo_2_4, p_wishbone_rx_fifo_fifo_2_5,
         p_wishbone_rx_fifo_fifo_2_6, p_wishbone_rx_fifo_fifo_2_7,
         p_wishbone_rx_fifo_fifo_2_8, p_wishbone_rx_fifo_fifo_2_9,
         p_wishbone_rx_fifo_fifo_2_10, p_wishbone_rx_fifo_fifo_2_11,
         p_wishbone_rx_fifo_fifo_2_12, p_wishbone_rx_fifo_fifo_2_13,
         p_wishbone_rx_fifo_fifo_2_14, p_wishbone_rx_fifo_fifo_2_15,
         p_wishbone_rx_fifo_fifo_2_16, p_wishbone_rx_fifo_fifo_2_17,
         p_wishbone_rx_fifo_fifo_2_18, p_wishbone_rx_fifo_fifo_2_19,
         p_wishbone_rx_fifo_fifo_2_20, p_wishbone_rx_fifo_fifo_2_21,
         p_wishbone_rx_fifo_fifo_2_22, p_wishbone_rx_fifo_fifo_2_23,
         p_wishbone_rx_fifo_fifo_2_24, p_wishbone_rx_fifo_fifo_2_25,
         p_wishbone_rx_fifo_fifo_2_26, p_wishbone_rx_fifo_fifo_2_27,
         p_wishbone_rx_fifo_fifo_2_28, p_wishbone_rx_fifo_fifo_2_29,
         p_wishbone_rx_fifo_fifo_2_30, p_wishbone_rx_fifo_fifo_2_31,
         p_wishbone_rx_fifo_fifo_1_0, p_wishbone_rx_fifo_fifo_1_1,
         p_wishbone_rx_fifo_fifo_1_2, p_wishbone_rx_fifo_fifo_1_3,
         p_wishbone_rx_fifo_fifo_1_4, p_wishbone_rx_fifo_fifo_1_5,
         p_wishbone_rx_fifo_fifo_1_6, p_wishbone_rx_fifo_fifo_1_7,
         p_wishbone_rx_fifo_fifo_1_8, p_wishbone_rx_fifo_fifo_1_9,
         p_wishbone_rx_fifo_fifo_1_10, p_wishbone_rx_fifo_fifo_1_11,
         p_wishbone_rx_fifo_fifo_1_12, p_wishbone_rx_fifo_fifo_1_13,
         p_wishbone_rx_fifo_fifo_1_14, p_wishbone_rx_fifo_fifo_1_15,
         p_wishbone_rx_fifo_fifo_1_16, p_wishbone_rx_fifo_fifo_1_17,
         p_wishbone_rx_fifo_fifo_1_18, p_wishbone_rx_fifo_fifo_1_19,
         p_wishbone_rx_fifo_fifo_1_20, p_wishbone_rx_fifo_fifo_1_21,
         p_wishbone_rx_fifo_fifo_1_22, p_wishbone_rx_fifo_fifo_1_23,
         p_wishbone_rx_fifo_fifo_1_24, p_wishbone_rx_fifo_fifo_1_25,
         p_wishbone_rx_fifo_fifo_1_26, p_wishbone_rx_fifo_fifo_1_27,
         p_wishbone_rx_fifo_fifo_1_28, p_wishbone_rx_fifo_fifo_1_29,
         p_wishbone_rx_fifo_fifo_1_30, p_wishbone_rx_fifo_fifo_1_31,
         p_wishbone_rx_fifo_fifo_0_0, p_wishbone_rx_fifo_fifo_0_1,
         p_wishbone_rx_fifo_fifo_0_2, p_wishbone_rx_fifo_fifo_0_3,
         p_wishbone_rx_fifo_fifo_0_4, p_wishbone_rx_fifo_fifo_0_5,
         p_wishbone_rx_fifo_fifo_0_6, p_wishbone_rx_fifo_fifo_0_7,
         p_wishbone_rx_fifo_fifo_0_8, p_wishbone_rx_fifo_fifo_0_9,
         p_wishbone_rx_fifo_fifo_0_10, p_wishbone_rx_fifo_fifo_0_11,
         p_wishbone_rx_fifo_fifo_0_12, p_wishbone_rx_fifo_fifo_0_13,
         p_wishbone_rx_fifo_fifo_0_14, p_wishbone_rx_fifo_fifo_0_15,
         p_wishbone_rx_fifo_fifo_0_16, p_wishbone_rx_fifo_fifo_0_17,
         p_wishbone_rx_fifo_fifo_0_18, p_wishbone_rx_fifo_fifo_0_19,
         p_wishbone_rx_fifo_fifo_0_20, p_wishbone_rx_fifo_fifo_0_21,
         p_wishbone_rx_fifo_fifo_0_22, p_wishbone_rx_fifo_fifo_0_23,
         p_wishbone_rx_fifo_fifo_0_24, p_wishbone_rx_fifo_fifo_0_25,
         p_wishbone_rx_fifo_fifo_0_26, p_wishbone_rx_fifo_fifo_0_27,
         p_wishbone_rx_fifo_fifo_0_28, p_wishbone_rx_fifo_fifo_0_29,
         p_wishbone_rx_fifo_fifo_0_30, p_wishbone_rx_fifo_fifo_0_31,
         p_wishbone_rx_fifo_write_pointer_3,
         p_wishbone_rx_fifo_write_pointer_2,
         p_wishbone_rx_fifo_write_pointer_1,
         p_wishbone_rx_fifo_write_pointer_0, p_wishbone_rx_fifo_N17,
         p_wishbone_rx_fifo_N16, p_wishbone_rx_fifo_N15,
         p_wishbone_rx_fifo_N14, p_wishbone_rxfifo_cnt_4,
         p_wishbone_rxfifo_cnt_3, p_wishbone_rxfifo_cnt_2,
         p_wishbone_rxfifo_cnt_1, p_wishbone_rxfifo_cnt_0;
  output wb_dat_o_0, wb_dat_o_1, wb_dat_o_2, wb_dat_o_3, wb_dat_o_4,
         wb_dat_o_5, wb_dat_o_6, wb_dat_o_7, wb_dat_o_8, wb_dat_o_9,
         wb_dat_o_10, wb_dat_o_11, wb_dat_o_12, wb_dat_o_13, wb_dat_o_14,
         wb_dat_o_15, wb_dat_o_16, wb_dat_o_17, wb_dat_o_18, wb_dat_o_19,
         wb_dat_o_20, wb_dat_o_21, wb_dat_o_22, wb_dat_o_23, wb_dat_o_24,
         wb_dat_o_25, wb_dat_o_26, wb_dat_o_27, wb_dat_o_28, wb_dat_o_29,
         wb_dat_o_30, wb_dat_o_31, m_wb_adr_o_0, m_wb_adr_o_1, m_wb_adr_o_2,
         m_wb_adr_o_3, m_wb_adr_o_4, m_wb_adr_o_5, m_wb_adr_o_6, m_wb_adr_o_7,
         m_wb_adr_o_8, m_wb_adr_o_9, m_wb_adr_o_10, m_wb_adr_o_11,
         m_wb_adr_o_12, m_wb_adr_o_13, m_wb_adr_o_14, m_wb_adr_o_15,
         m_wb_adr_o_16, m_wb_adr_o_17, m_wb_adr_o_18, m_wb_adr_o_19,
         m_wb_adr_o_20, m_wb_adr_o_21, m_wb_adr_o_22, m_wb_adr_o_23,
         m_wb_adr_o_24, m_wb_adr_o_25, m_wb_adr_o_26, m_wb_adr_o_27,
         m_wb_adr_o_28, m_wb_adr_o_29, m_wb_adr_o_30, m_wb_adr_o_31,
         m_wb_sel_o_0, m_wb_sel_o_1, m_wb_sel_o_2, m_wb_sel_o_3, m_wb_dat_o_0,
         m_wb_dat_o_1, m_wb_dat_o_2, m_wb_dat_o_3, m_wb_dat_o_4, m_wb_dat_o_5,
         m_wb_dat_o_6, m_wb_dat_o_7, m_wb_dat_o_8, m_wb_dat_o_9, m_wb_dat_o_10,
         m_wb_dat_o_11, m_wb_dat_o_12, m_wb_dat_o_13, m_wb_dat_o_14,
         m_wb_dat_o_15, m_wb_dat_o_16, m_wb_dat_o_17, m_wb_dat_o_18,
         m_wb_dat_o_19, m_wb_dat_o_20, m_wb_dat_o_21, m_wb_dat_o_22,
         m_wb_dat_o_23, m_wb_dat_o_24, m_wb_dat_o_25, m_wb_dat_o_26,
         m_wb_dat_o_27, m_wb_dat_o_28, m_wb_dat_o_29, m_wb_dat_o_30,
         m_wb_dat_o_31, mtxd_pad_o_0, mtxd_pad_o_1, mtxd_pad_o_2, mtxd_pad_o_3,
         wb_ack_o, wb_err_o, m_wb_we_o, m_wb_cyc_o, m_wb_stb_o, mtxen_pad_o,
         mtxerr_pad_o, mdc_pad_o, md_pad_o, md_padoe_o, int_o, N10,
         RxAbortRst_sync1, n126, WillSendControlFrame, N23, N24, N25, n124,
         n125, WillTransmit, N9, temp_wb_dat_o_0, temp_wb_dat_o_1,
         temp_wb_dat_o_2, temp_wb_dat_o_3, temp_wb_dat_o_4, temp_wb_dat_o_5,
         temp_wb_dat_o_6, temp_wb_dat_o_7, temp_wb_dat_o_8, temp_wb_dat_o_9,
         temp_wb_dat_o_10, temp_wb_dat_o_11, temp_wb_dat_o_12,
         temp_wb_dat_o_13, temp_wb_dat_o_14, temp_wb_dat_o_15,
         temp_wb_dat_o_16, temp_wb_dat_o_17, temp_wb_dat_o_18,
         temp_wb_dat_o_19, temp_wb_dat_o_20, temp_wb_dat_o_21,
         temp_wb_dat_o_22, temp_wb_dat_o_23, temp_wb_dat_o_24,
         temp_wb_dat_o_25, temp_wb_dat_o_26, temp_wb_dat_o_27,
         temp_wb_dat_o_28, temp_wb_dat_o_29, temp_wb_dat_o_30,
         temp_wb_dat_o_31, p_miim1_n133, p_miim1_n134, p_miim1_n135,
         p_miim1_n136, p_miim1_n153, p_miim1_n137, p_miim1_n138, p_miim1_n139,
         p_miim1_n140, p_miim1_n141, p_miim1_n142, p_miim1_n156, p_miim1_N9,
         p_miim1_n143, p_miim1_n144, p_miim1_n145, p_miim1_n154, p_miim1_n146,
         p_miim1_n147, p_miim1_n155, p_miim1_EndBusy_d, p_miim1_N8,
         p_miim1_n148, p_miim1_n149, p_miim1_n150, p_miim1_n157, p_miim1_n151,
         p_miim1_WCtrlData_q2, p_miim1_WCtrlData_q1, r_WCtrlData,
         p_miim1_RStat_q2, p_miim1_RStat_q1, r_RStat, p_miim1_n152,
         p_miim1_ScanStat_q1, r_ScanStat, p_ethreg1_n678, p_ethreg1_n679,
         p_ethreg1_n680, p_ethreg1_n681, p_ethreg1_n682, p_ethreg1_n683,
         p_ethreg1_n684, p_ethreg1_N228, p_ethreg1_ResetRxCIrq_sync1,
         p_ethreg1_SetRxCIrq_sync2, p_ethreg1_SetRxCIrq_sync1,
         p_ethreg1_SetRxCIrq_rxclk, p_ethreg1_n685, p_ethreg1_N222,
         p_ethreg1_SetTxCIrq_sync2, p_ethreg1_SetTxCIrq_sync1,
         p_ethreg1_SetTxCIrq_txclk, p_ethreg1_n686, p_maccontrol1_n53,
         p_maccontrol1_n54, TxDoneIn, TxAbortIn, p_maccontrol1_n55,
         p_txethmac1_n152, p_txethmac1_n153, p_txethmac1_n149,
         p_txethmac1_PacketFinished_d, p_txethmac1_n148, p_txethmac1_n147,
         p_txethmac1_n150, p_txethmac1_n155, p_txethmac1_MTxD_d_0,
         p_txethmac1_MTxD_d_1, p_txethmac1_MTxD_d_2, p_txethmac1_MTxD_d_3,
         p_txethmac1_N88, p_txethmac1_N86, p_txethmac1_N87, p_txethmac1_n156,
         p_txethmac1_N29, p_txethmac1_n151, p_txethmac1_n154, p_rxethmac1_n95,
         p_rxethmac1_n94, p_rxethmac1_N51, p_rxethmac1_GenerateRxEndFrm,
         p_rxethmac1_RxStartFrm_d, p_rxethmac1_GenerateRxStartFrm,
         p_rxethmac1_RxValid_d, n33940, p_rxethmac1_RxData_d_7,
         p_rxethmac1_n103, p_rxethmac1_RxData_d_6, p_rxethmac1_n102,
         p_rxethmac1_RxData_d_5, p_rxethmac1_n101, p_rxethmac1_RxData_d_4,
         p_rxethmac1_n100, p_rxethmac1_RxData_d_3, p_rxethmac1_n99,
         p_rxethmac1_RxData_d_2, p_rxethmac1_n98, p_rxethmac1_RxData_d_1,
         p_rxethmac1_n97, p_rxethmac1_RxData_d_0, p_rxethmac1_n96,
         RxStateData_0, p_rxethmac1_LatchedByte_4, p_rxethmac1_LatchedByte_5,
         p_rxethmac1_LatchedByte_6, p_rxethmac1_LatchedByte_7, MRxD_Lb_0,
         MRxD_Lb_1, MRxD_Lb_2, MRxD_Lb_3, p_rxethmac1_n104, p_rxethmac1_n105,
         p_rxethmac1_n106, p_rxethmac1_n107, p_rxethmac1_n108,
         p_rxethmac1_n109, p_rxethmac1_N3, p_wishbone_Busy_IRQ_sync2,
         p_wishbone_Busy_IRQ_sync1, p_wishbone_Busy_IRQ_rck, p_wishbone_n2138,
         p_wishbone_N1329, p_wishbone_N1326, p_wishbone_N1322,
         p_wishbone_N1319, RxStatusWriteLatched_sync2,
         p_wishbone_RxStatusWriteLatched_sync1,
         p_wishbone_RxStatusWriteLatched, p_wishbone_n2139, p_wishbone_n2141,
         p_wishbone_n2142, p_wishbone_n2143, p_wishbone_n2144,
         p_wishbone_n2145, p_wishbone_n2146, p_wishbone_n2147,
         p_wishbone_n2148, p_wishbone_n2149, p_wishbone_n2150,
         p_wishbone_n2151, p_wishbone_n2152, p_wishbone_n2153,
         p_wishbone_n2154, p_wishbone_n2155, p_wishbone_n2156,
         p_wishbone_n2157, p_wishbone_n2158, p_wishbone_n2159,
         p_wishbone_n2160, p_wishbone_n2161, p_wishbone_n2162,
         p_wishbone_n2163, p_wishbone_n2164, p_wishbone_n2165,
         p_wishbone_n2166, p_wishbone_n2167, p_wishbone_n2168,
         p_wishbone_n2169, p_wishbone_n2140, p_wishbone_n2171,
         p_wishbone_n2172, p_wishbone_n2173, p_wishbone_n2174,
         p_wishbone_n2175, p_wishbone_n2176, p_wishbone_n2177,
         p_wishbone_n2178, p_wishbone_n2179, p_wishbone_n2180,
         p_wishbone_n2181, p_wishbone_n2182, p_wishbone_n2183,
         p_wishbone_n2184, p_wishbone_n2185, p_wishbone_n2186,
         p_wishbone_n2187, p_wishbone_n2188, p_wishbone_n2189,
         p_wishbone_n2190, p_wishbone_n2191, p_wishbone_n2192,
         p_wishbone_n2193, p_wishbone_n2194, p_wishbone_n2195,
         p_wishbone_n2196, p_wishbone_n2197, p_wishbone_n2198,
         p_wishbone_n2199, p_wishbone_n2170, p_wishbone_n2201,
         p_wishbone_n2202, p_wishbone_n2203, p_wishbone_n2204,
         p_wishbone_n2205, p_wishbone_n2206, p_wishbone_n2207,
         p_wishbone_n2208, p_wishbone_n2209, p_wishbone_n2210,
         p_wishbone_n2211, p_wishbone_n2212, p_wishbone_n2213,
         p_wishbone_n2214, p_wishbone_n2215, p_wishbone_n2216,
         p_wishbone_n2217, p_wishbone_n2218, p_wishbone_n2219,
         p_wishbone_n2220, p_wishbone_n2221, p_wishbone_n2222,
         p_wishbone_n2223, p_wishbone_n2224, p_wishbone_n2225,
         p_wishbone_n2226, p_wishbone_n2227, p_wishbone_n2228,
         p_wishbone_n2229, p_wishbone_n2200, p_wishbone_n2339,
         p_wishbone_n2333, p_wishbone_n2334, p_wishbone_n2342,
         p_wishbone_n2341, p_wishbone_n2335, p_wishbone_n2336,
         p_wishbone_n2337, p_wishbone_n2340, p_wishbone_n2462,
         p_wishbone_n2250, p_wishbone_n2258, p_wishbone_n2251,
         p_wishbone_n2259, p_wishbone_n2252, p_wishbone_n2260,
         p_wishbone_n2253, p_wishbone_n2261, p_wishbone_n2254,
         p_wishbone_n2262, p_wishbone_n2255, p_wishbone_n2263,
         p_wishbone_n2256, p_wishbone_n2264, p_wishbone_n2257,
         p_wishbone_n2265, p_wishbone_n2266, p_wishbone_n2267,
         p_wishbone_n2268, p_wishbone_n2269, p_wishbone_n2270,
         p_wishbone_n2271, p_wishbone_n2272, p_wishbone_n2273,
         p_wishbone_n2274, p_wishbone_n2275, p_wishbone_n2276,
         p_wishbone_n2277, p_wishbone_n2278, p_wishbone_n2279,
         p_wishbone_n2280, p_wishbone_n2281, p_wishbone_n2282,
         p_wishbone_n2283, p_wishbone_n2284, p_wishbone_n2285,
         p_wishbone_n2286, p_wishbone_n2287, p_wishbone_n2288,
         p_wishbone_n2289, p_wishbone_n2290, p_wishbone_n2291,
         p_wishbone_n2292, p_wishbone_n2293, p_wishbone_TxStartFrm_syncb1,
         p_wishbone_TxStartFrm_sync2, p_wishbone_TxStartFrm_sync1,
         p_wishbone_TxStartFrm_wb, p_wishbone_n2294, p_wishbone_n2295,
         p_wishbone_n2437, p_wishbone_n2230, p_wishbone_n2231,
         p_wishbone_n2249, n33933, p_wishbone_BlockingTxStatusWrite_sync2,
         p_wishbone_BlockingTxStatusWrite_sync1,
         p_wishbone_BlockingTxStatusWrite, p_wishbone_n2232, p_wishbone_n2239,
         p_wishbone_n2233, p_wishbone_n2241, p_wishbone_n2234,
         p_wishbone_n2242, p_wishbone_n2235, p_wishbone_n2243,
         p_wishbone_n2236, p_wishbone_n2244, p_wishbone_n2237,
         p_wishbone_n2245, p_wishbone_n2238, p_wishbone_n2246,
         p_wishbone_n2247, p_wishbone_n2347, p_wishbone_n2240,
         p_wishbone_n2085, p_wishbone_n2086, p_wishbone_n2441,
         p_wishbone_n2327, p_wishbone_n2328, p_wishbone_n2329, p_wishbone_N75,
         p_wishbone_n2331, p_wishbone_n2469, p_wishbone_n2456,
         p_wishbone_n2455, p_wishbone_n2454, p_wishbone_n2453,
         p_wishbone_n2452, p_wishbone_n2451, p_wishbone_n2450,
         p_wishbone_n2449, p_wishbone_n2448, p_wishbone_n2447,
         p_wishbone_n2446, p_wishbone_n2445, p_wishbone_n2444,
         p_wishbone_n2443, p_wishbone_n2442, p_wishbone_n2440,
         p_wishbone_n2439, p_wishbone_n2438, p_wishbone_n2436,
         p_wishbone_n2434, p_wishbone_n2433, p_wishbone_n2432,
         p_wishbone_n2431, p_wishbone_n2430, p_wishbone_n2429,
         p_wishbone_n2324, p_wishbone_n2323, p_wishbone_n2322,
         p_wishbone_n2321, p_wishbone_n2087, p_wishbone_n2418,
         p_wishbone_n2419, p_wishbone_n2420, p_wishbone_n2421,
         p_wishbone_n2422, p_wishbone_n2423, p_wishbone_n2424,
         p_wishbone_n2088, p_wishbone_n2325, p_wishbone_n2382,
         p_wishbone_n2406, p_wishbone_n2381, p_wishbone_n2405,
         p_wishbone_n2380, p_wishbone_n2404, p_wishbone_n2379,
         p_wishbone_n2403, p_wishbone_n2378, p_wishbone_n2402,
         p_wishbone_n2377, p_wishbone_n2401, p_wishbone_n2376,
         p_wishbone_n2400, p_wishbone_n2375, p_wishbone_n2399,
         p_wishbone_n2365, p_wishbone_n2366, p_wishbone_n2363,
         p_wishbone_n2364, p_wishbone_n2361, p_wishbone_n2362,
         p_wishbone_n2359, p_wishbone_n2360, p_wishbone_n2357,
         p_wishbone_n2358, p_wishbone_n2355, p_wishbone_n2356,
         p_wishbone_n2353, p_wishbone_n2354, p_wishbone_n2351,
         p_wishbone_n2352, p_wishbone_n2373, p_wishbone_n2372,
         p_wishbone_n2371, p_wishbone_n2370, p_wishbone_n2369,
         p_wishbone_n2368, p_wishbone_n2367, p_wishbone_n2390,
         p_wishbone_n2389, p_wishbone_n2388, p_wishbone_n2387,
         p_wishbone_n2386, p_wishbone_n2385, p_wishbone_n2384,
         p_wishbone_n2383, p_wishbone_WriteRxDataToFifoSync2,
         p_wishbone_WriteRxDataToFifoSync1, p_wishbone_WriteRxDataToFifo,
         p_wishbone_n2413, p_wishbone_n2414, p_wishbone_n2411,
         p_wishbone_n2410, p_wishbone_ShiftEndedSync_c1,
         p_wishbone_ShiftEndedSync2, p_wishbone_ShiftEndedSync1,
         p_wishbone_ShiftEnded_rck, p_wishbone_n2412, p_wishbone_n2407,
         p_wishbone_n2408, p_wishbone_n2409, p_wishbone_n2425,
         p_wishbone_n2426, p_wishbone_n2427, p_wishbone_n2374,
         p_wishbone_n2398, p_wishbone_n2397, p_wishbone_n2396,
         p_wishbone_n2395, p_wishbone_n2394, p_wishbone_n2393,
         p_wishbone_n2392, p_wishbone_n2391, p_wishbone_n2416,
         p_wishbone_n2415, p_wishbone_n2417, p_wishbone_n2326, p_wishbone_RxEn,
         p_wishbone_n2428, p_wishbone_n2332, p_wishbone_WbEn, p_wishbone_n2330,
         p_wishbone_n2089, p_wishbone_n2090, p_wishbone_n2091,
         p_wishbone_n2092, p_wishbone_n2093, p_wishbone_n2094,
         p_wishbone_n2095, p_wishbone_n2096, p_wishbone_n2097,
         p_wishbone_n2098, p_wishbone_n2099, p_wishbone_n2100,
         p_wishbone_n2101, p_wishbone_n2102, p_wishbone_n2103,
         p_wishbone_n2104, p_wishbone_n2248, p_wishbone_n2320,
         p_wishbone_n2301, p_wishbone_n2302, p_wishbone_n2303,
         p_wishbone_n2304, p_wishbone_n2305, p_wishbone_n2306,
         p_wishbone_n2307, p_wishbone_n2308, p_wishbone_n2309,
         p_wishbone_n2310, p_wishbone_n2311, p_wishbone_n2312,
         p_wishbone_n2313, p_wishbone_n2314, p_wishbone_n2299,
         p_wishbone_n2315, p_wishbone_n2316, p_wishbone_n2105,
         p_wishbone_n2106, p_wishbone_n2107, p_wishbone_n2108,
         p_wishbone_n2319, p_wishbone_TxEn, p_wishbone_n2457, p_wishbone_n2458,
         p_wishbone_n2318, p_wishbone_n2317, p_wishbone_n2459,
         p_wishbone_n2460, p_wishbone_n2461, p_wishbone_n2348, p_wishbone_N867,
         p_wishbone_n2349, n33934, p_wishbone_n2463, p_wishbone_n2343,
         p_wishbone_n2344, p_wishbone_n2345, p_wishbone_n2346,
         p_wishbone_n2350, p_wishbone_n2466, p_wishbone_n2338,
         p_wishbone_n2464, p_wishbone_n2465, p_wishbone_n2467,
         p_wishbone_ReadTxDataFromFifo_sync2,
         p_wishbone_ReadTxDataFromFifo_syncb2,
         p_wishbone_ReadTxDataFromFifo_syncb1,
         p_wishbone_ReadTxDataFromFifo_sync1,
         p_wishbone_ReadTxDataFromFifo_tck, p_wishbone_n2296, p_wishbone_n2297,
         p_wishbone_n2298, p_wishbone_n2300, p_wishbone_LatchValidBytes,
         p_wishbone_N811, p_wishbone_n2468, p_wishbone_n2435, p_wishbone_n2109,
         p_wishbone_n2470, p_wishbone_n2110, p_wishbone_n2111,
         p_wishbone_n2112, p_wishbone_n2113, p_wishbone_n2114,
         p_wishbone_n2115, p_wishbone_n2116, p_wishbone_n2117,
         p_wishbone_n2118, p_wishbone_n2119, p_wishbone_n2120,
         p_wishbone_n2121, p_wishbone_n2122, p_wishbone_n2123,
         p_wishbone_n2124, p_wishbone_n2125, p_wishbone_n2126,
         p_wishbone_n2127, p_wishbone_n2128, p_wishbone_n2129,
         p_wishbone_n2130, p_wishbone_n2131, p_wishbone_n2132,
         p_wishbone_n2133, p_wishbone_RxAbortSyncb1, p_wishbone_RxAbortSync2,
         p_wishbone_RxAbortSync3, p_wishbone_RxAbortSync1,
         p_wishbone_RxAbortLatched, p_wishbone_n2471, p_wishbone_n2472,
         p_wishbone_SyncRxStartFrm_q, p_wishbone_LatchedRxStartFrm,
         p_wishbone_n2473, p_wishbone_TxAbort_wb, p_wishbone_TxAbortSync1,
         TxAbort, p_wishbone_TxDone_wb, p_wishbone_TxDoneSync1, TxDone,
         p_wishbone_TxRetry_wb, p_wishbone_TxRetrySync1, n33935,
         p_wishbone_n2474, r_RxEn, r_TxEn, p_macstatus1_n89, p_macstatus1_n90,
         p_macstatus1_n82, p_macstatus1_n83, p_macstatus1_n84,
         p_macstatus1_n85, p_macstatus1_n86, p_macstatus1_n87,
         p_macstatus1_n91, p_macstatus1_n92, p_macstatus1_n93,
         p_macstatus1_n94, p_macstatus1_n95, p_macstatus1_n96, LoadRxStatus,
         p_macstatus1_TakeSample, p_macstatus1_N7, p_macstatus1_n97,
         p_miim1_clkgen_n35, p_miim1_clkgen_N21, p_miim1_clkgen_N20,
         p_miim1_clkgen_N19, p_miim1_clkgen_N18, p_miim1_clkgen_N17,
         p_miim1_clkgen_N16, p_miim1_clkgen_N15, p_miim1_shftrg_n145,
         p_miim1_shftrg_n146, p_miim1_shftrg_n147, p_miim1_shftrg_n148,
         p_miim1_shftrg_n149, p_miim1_shftrg_n150, p_miim1_shftrg_n151,
         p_miim1_shftrg_n152, p_miim1_shftrg_n153, p_miim1_shftrg_n154,
         p_miim1_shftrg_n155, p_miim1_shftrg_n156, p_miim1_shftrg_n157,
         p_miim1_shftrg_n158, p_miim1_shftrg_n159, p_miim1_shftrg_n160,
         p_miim1_shftrg_n161, p_miim1_shftrg_n137, p_miim1_shftrg_n138,
         p_miim1_shftrg_n139, p_miim1_shftrg_n140, p_miim1_shftrg_n141,
         p_miim1_shftrg_n142, p_miim1_shftrg_n143, p_miim1_shftrg_n144,
         p_miim1_outctrl_n33, p_miim1_outctrl_n34, p_miim1_outctrl_n35,
         p_miim1_outctrl_n36, p_miim1_outctrl_n37, p_miim1_outctrl_n38,
         p_ethreg1_MODER_0_n21, p_ethreg1_MODER_0_n22, p_ethreg1_MODER_0_n23,
         p_ethreg1_MODER_0_n24, p_ethreg1_MODER_0_n25, p_ethreg1_MODER_0_n26,
         p_ethreg1_MODER_0_n27, p_ethreg1_MODER_0_n28, p_ethreg1_MODER_1_n23,
         p_ethreg1_MODER_1_n24, p_ethreg1_MODER_1_n25, p_ethreg1_MODER_1_n26,
         p_ethreg1_MODER_1_n27, n33922, p_ethreg1_MODER_1_n29, n33921, n33920,
         p_ethreg1_INT_MASK_0_n19, p_ethreg1_INT_MASK_0_n20,
         p_ethreg1_INT_MASK_0_n21, p_ethreg1_INT_MASK_0_n22,
         p_ethreg1_INT_MASK_0_n23, p_ethreg1_INT_MASK_0_n24,
         p_ethreg1_INT_MASK_0_n25, p_ethreg1_IPGT_0_n21, n33931,
         p_ethreg1_IPGT_0_n23, p_ethreg1_IPGT_0_n24, n33927,
         p_ethreg1_IPGT_0_n26, p_ethreg1_IPGT_0_n27, p_ethreg1_IPGR1_0_n21,
         p_ethreg1_IPGR1_0_n22, n33929, n33928, p_ethreg1_IPGR1_0_n25,
         p_ethreg1_IPGR1_0_n26, p_ethreg1_IPGR1_0_n27,
         p_ethreg1_PACKETLEN_1_n23, n33924, n33923, p_ethreg1_PACKETLEN_1_n26,
         p_ethreg1_PACKETLEN_1_n27, p_ethreg1_PACKETLEN_1_n28,
         p_ethreg1_PACKETLEN_1_n29, p_ethreg1_PACKETLEN_1_n30,
         p_ethreg1_PACKETLEN_2_n22, p_ethreg1_PACKETLEN_2_n23,
         p_ethreg1_PACKETLEN_2_n24, p_ethreg1_PACKETLEN_2_n25,
         p_ethreg1_PACKETLEN_2_n26, p_ethreg1_PACKETLEN_2_n27,
         p_ethreg1_PACKETLEN_2_n17, p_ethreg1_PACKETLEN_2_n29,
         p_ethreg1_COLLCONF_0_n21, p_ethreg1_COLLCONF_0_n22,
         p_ethreg1_COLLCONF_0_n23, p_ethreg1_COLLCONF_0_n24,
         p_ethreg1_COLLCONF_0_n25, p_ethreg1_COLLCONF_0_n26,
         p_ethreg1_COLLCONF_2_n15, p_ethreg1_COLLCONF_2_n16,
         p_ethreg1_COLLCONF_2_n17, p_ethreg1_COLLCONF_2_n18,
         p_ethreg1_CTRLMODER_0_n10, p_ethreg1_CTRLMODER_0_n11,
         p_ethreg1_CTRLMODER_0_n12, p_ethreg1_MIIMODER_0_n24,
         p_ethreg1_MIIMODER_0_n25, p_ethreg1_MIIMODER_0_n26,
         p_ethreg1_MIIMODER_0_n27, p_ethreg1_MIIMODER_0_n28,
         p_ethreg1_MIIMODER_0_n29, p_ethreg1_MIIMODER_0_n30,
         p_ethreg1_MIIMODER_0_n31, n33932, p_ethreg1_MIIADDRESS_0_n15,
         p_ethreg1_MIIADDRESS_0_n16, p_ethreg1_MIIADDRESS_0_n17,
         p_ethreg1_MIIADDRESS_0_n18, p_ethreg1_MIIADDRESS_0_n19,
         p_ethreg1_MIIRX_DATA_n37, p_ethreg1_MIIRX_DATA_n38,
         p_ethreg1_MIIRX_DATA_n39, p_ethreg1_MIIRX_DATA_n40,
         p_ethreg1_MIIRX_DATA_n41, p_ethreg1_MIIRX_DATA_n42,
         p_ethreg1_MIIRX_DATA_n43, p_ethreg1_MIIRX_DATA_n44,
         p_ethreg1_MIIRX_DATA_n45, p_ethreg1_MIIRX_DATA_n46,
         p_ethreg1_MIIRX_DATA_n47, p_ethreg1_MIIRX_DATA_n48,
         p_ethreg1_MIIRX_DATA_n49, p_ethreg1_MIIRX_DATA_n50,
         p_ethreg1_MIIRX_DATA_n51, p_ethreg1_MIIRX_DATA_n52,
         p_maccontrol1_receivecontrol1_n503,
         p_maccontrol1_receivecontrol1_n507,
         p_maccontrol1_receivecontrol1_n506,
         p_maccontrol1_receivecontrol1_n505,
         p_maccontrol1_receivecontrol1_n504,
         p_maccontrol1_receivecontrol1_n524,
         p_maccontrol1_receivecontrol1_n501,
         p_maccontrol1_receivecontrol1_PauseTimerEq0_sync1, n33939,
         p_maccontrol1_receivecontrol1_N208,
         p_maccontrol1_receivecontrol1_n508,
         p_maccontrol1_receivecontrol1_n509,
         p_maccontrol1_receivecontrol1_n510,
         p_maccontrol1_receivecontrol1_n511,
         p_maccontrol1_receivecontrol1_n512,
         p_maccontrol1_receivecontrol1_n513,
         p_maccontrol1_receivecontrol1_n514,
         p_maccontrol1_receivecontrol1_n515,
         p_maccontrol1_receivecontrol1_n516,
         p_maccontrol1_receivecontrol1_n517,
         p_maccontrol1_receivecontrol1_n518,
         p_maccontrol1_receivecontrol1_n519,
         p_maccontrol1_receivecontrol1_n520,
         p_maccontrol1_receivecontrol1_n521,
         p_maccontrol1_receivecontrol1_n522,
         p_maccontrol1_receivecontrol1_n523,
         p_maccontrol1_receivecontrol1_n525,
         p_maccontrol1_receivecontrol1_n541,
         p_maccontrol1_receivecontrol1_n540,
         p_maccontrol1_receivecontrol1_n539,
         p_maccontrol1_receivecontrol1_n538,
         p_maccontrol1_receivecontrol1_n537,
         p_maccontrol1_receivecontrol1_n536,
         p_maccontrol1_receivecontrol1_n535,
         p_maccontrol1_receivecontrol1_n534,
         p_maccontrol1_receivecontrol1_n533,
         p_maccontrol1_receivecontrol1_n532,
         p_maccontrol1_receivecontrol1_n531,
         p_maccontrol1_receivecontrol1_n530,
         p_maccontrol1_receivecontrol1_n529,
         p_maccontrol1_receivecontrol1_n528,
         p_maccontrol1_receivecontrol1_n527,
         p_maccontrol1_receivecontrol1_n526,
         p_maccontrol1_receivecontrol1_n558,
         p_maccontrol1_receivecontrol1_n559,
         p_maccontrol1_receivecontrol1_n561,
         p_maccontrol1_receivecontrol1_n560,
         p_maccontrol1_receivecontrol1_n557,
         p_maccontrol1_receivecontrol1_n556,
         p_maccontrol1_receivecontrol1_n555,
         p_maccontrol1_receivecontrol1_n554,
         p_maccontrol1_receivecontrol1_n553,
         p_maccontrol1_receivecontrol1_n552,
         p_maccontrol1_receivecontrol1_n551,
         p_maccontrol1_receivecontrol1_n550,
         p_maccontrol1_receivecontrol1_n549,
         p_maccontrol1_receivecontrol1_n548,
         p_maccontrol1_receivecontrol1_n547,
         p_maccontrol1_receivecontrol1_n546,
         p_maccontrol1_receivecontrol1_n545,
         p_maccontrol1_receivecontrol1_n544,
         p_maccontrol1_receivecontrol1_n543,
         p_maccontrol1_receivecontrol1_n542,
         p_maccontrol1_receivecontrol1_n564,
         p_maccontrol1_receivecontrol1_n563,
         p_maccontrol1_receivecontrol1_n562,
         p_maccontrol1_receivecontrol1_n566,
         p_maccontrol1_receivecontrol1_n565,
         p_maccontrol1_receivecontrol1_n567,
         p_maccontrol1_receivecontrol1_n568,
         p_maccontrol1_receivecontrol1_n569,
         p_maccontrol1_receivecontrol1_n570,
         p_maccontrol1_transmitcontrol1_n263,
         p_maccontrol1_transmitcontrol1_n264,
         p_maccontrol1_transmitcontrol1_n265,
         p_maccontrol1_transmitcontrol1_n266,
         p_maccontrol1_transmitcontrol1_n267,
         p_maccontrol1_transmitcontrol1_n268,
         p_maccontrol1_transmitcontrol1_n269,
         p_maccontrol1_transmitcontrol1_n270,
         p_maccontrol1_transmitcontrol1_n275,
         p_maccontrol1_transmitcontrol1_n274,
         p_maccontrol1_transmitcontrol1_n273,
         p_maccontrol1_transmitcontrol1_n272,
         p_maccontrol1_transmitcontrol1_n283,
         p_maccontrol1_transmitcontrol1_n276,
         p_maccontrol1_transmitcontrol1_n277,
         p_maccontrol1_transmitcontrol1_n278,
         p_maccontrol1_transmitcontrol1_n279,
         p_maccontrol1_transmitcontrol1_n271, p_maccontrol1_TxCtrlStartFrm,
         p_maccontrol1_transmitcontrol1_n280,
         p_maccontrol1_transmitcontrol1_n281,
         p_maccontrol1_transmitcontrol1_n282,
         p_maccontrol1_transmitcontrol1_N31,
         p_maccontrol1_transmitcontrol1_n285,
         p_maccontrol1_transmitcontrol1_n284, p_txethmac1_txcounters1_n172,
         p_txethmac1_txcounters1_n173, p_txethmac1_txcounters1_n174,
         p_txethmac1_txcounters1_n188, p_txethmac1_txcounters1_n187,
         p_txethmac1_txcounters1_n186, p_txethmac1_txcounters1_n185,
         p_txethmac1_txcounters1_n184, p_txethmac1_txcounters1_n183,
         p_txethmac1_txcounters1_n182, p_txethmac1_txcounters1_n181,
         p_txethmac1_txcounters1_n180, p_txethmac1_txcounters1_n179,
         p_txethmac1_txcounters1_n178, p_txethmac1_txcounters1_n177,
         p_txethmac1_txcounters1_n176, p_txethmac1_txcounters1_n175,
         p_txethmac1_txcounters1_n189, p_txethmac1_txcounters1_n190,
         p_txethmac1_txcounters1_n191, p_txethmac1_txcounters1_n192,
         p_txethmac1_txcounters1_n193, p_txethmac1_txcounters1_n194,
         p_txethmac1_txcounters1_n195, p_txethmac1_txcounters1_n196,
         p_txethmac1_txcounters1_n197, p_txethmac1_txcounters1_n198,
         p_txethmac1_txcounters1_n199, p_txethmac1_txcounters1_n200,
         p_txethmac1_txcounters1_n201, p_txethmac1_txcounters1_n202,
         p_txethmac1_txcounters1_n204, p_txethmac1_txcounters1_n203,
         p_txethmac1_txcounters1_n205, p_txethmac1_txcounters1_n206,
         p_txethmac1_txstatem1_n90, p_txethmac1_StateJam,
         p_txethmac1_txstatem1_n93, p_txethmac1_txstatem1_n94,
         p_txethmac1_StartData_1, p_txethmac1_StartData_0,
         p_txethmac1_txstatem1_n95, p_txethmac1_txstatem1_n96,
         p_txethmac1_txstatem1_n97, p_txethmac1_txstatem1_n92,
         p_txethmac1_txstatem1_n91, p_txethmac1_txstatem1_n98,
         p_txethmac1_txcrc_N25, p_txethmac1_txcrc_N21, p_txethmac1_txcrc_N17,
         p_txethmac1_txcrc_N13, p_txethmac1_txcrc_N9, p_txethmac1_txcrc_N5,
         p_txethmac1_txcrc_N8, p_txethmac1_txcrc_N26, p_txethmac1_txcrc_N22,
         p_txethmac1_txcrc_N18, p_txethmac1_txcrc_N14, p_txethmac1_txcrc_N10,
         p_txethmac1_txcrc_N6, p_txethmac1_txcrc_N34, p_txethmac1_txcrc_N30,
         p_txethmac1_txcrc_N4, p_txethmac1_txcrc_N32, p_txethmac1_txcrc_N28,
         p_txethmac1_txcrc_N24, p_txethmac1_txcrc_N20, p_txethmac1_txcrc_N16,
         p_txethmac1_txcrc_N12, p_txethmac1_txcrc_N33, p_txethmac1_txcrc_N29,
         p_txethmac1_txcrc_N31, p_txethmac1_txcrc_N27, p_txethmac1_txcrc_N23,
         p_txethmac1_txcrc_N19, p_txethmac1_txcrc_N15, p_txethmac1_txcrc_N11,
         p_txethmac1_txcrc_N7, p_txethmac1_txcrc_N3, p_txethmac1_random1_n98,
         p_txethmac1_random1_n99, p_txethmac1_random1_n100,
         p_txethmac1_random1_n101, p_txethmac1_random1_n102,
         p_txethmac1_random1_n103, p_txethmac1_random1_n104,
         p_txethmac1_random1_n105, p_txethmac1_random1_n106,
         p_txethmac1_random1_n107, p_txethmac1_random1_x_8,
         p_txethmac1_random1_x_7, p_txethmac1_random1_x_6,
         p_txethmac1_random1_x_5, p_txethmac1_random1_x_4,
         p_txethmac1_random1_x_3, p_txethmac1_random1_x_2,
         p_txethmac1_random1_x_1, p_txethmac1_random1_x_0,
         p_txethmac1_random1_n108, p_rxethmac1_rxstatem1_n38,
         p_rxethmac1_rxstatem1_n37, p_rxethmac1_rxstatem1_n39,
         p_rxethmac1_rxstatem1_n40, p_rxethmac1_rxstatem1_n41,
         p_rxethmac1_rxstatem1_n42, p_rxethmac1_rxcounters1_n175,
         p_rxethmac1_rxcounters1_n174, p_rxethmac1_rxcounters1_n173,
         p_rxethmac1_rxcounters1_n172, p_rxethmac1_rxcounters1_n171,
         p_rxethmac1_rxcounters1_n170, p_rxethmac1_rxcounters1_n169,
         p_rxethmac1_rxcounters1_n168, p_rxethmac1_rxcounters1_n167,
         p_rxethmac1_rxcounters1_n166, p_rxethmac1_rxcounters1_n165,
         p_rxethmac1_rxcounters1_n164, p_rxethmac1_rxcounters1_n163,
         p_rxethmac1_rxcounters1_n162, p_rxethmac1_rxcounters1_n176,
         p_rxethmac1_rxcounters1_n161, p_rxethmac1_rxcounters1_n178,
         p_rxethmac1_rxcounters1_n177, p_rxethmac1_rxcounters1_n179,
         p_rxethmac1_rxcounters1_n180, p_rxethmac1_rxcounters1_n183,
         p_rxethmac1_rxcounters1_n182, p_rxethmac1_rxcounters1_n181,
         p_rxethmac1_rxcounters1_n184, p_rxethmac1_rxcounters1_n185,
         p_rxethmac1_rxaddrcheck1_n290, p_rxethmac1_rxaddrcheck1_n294,
         p_rxethmac1_rxaddrcheck1_N10, p_rxethmac1_rxaddrcheck1_n295,
         p_wishbone_bd_ram_n17793, p_wishbone_bd_ram_n17794,
         p_wishbone_bd_ram_n17795, p_wishbone_bd_ram_n17796,
         p_wishbone_bd_ram_n17797, p_wishbone_bd_ram_n17798,
         p_wishbone_bd_ram_n17799, p_wishbone_bd_ram_n17800,
         p_wishbone_bd_ram_n17801, p_wishbone_bd_ram_n17802,
         p_wishbone_bd_ram_n17803, p_wishbone_bd_ram_n17804,
         p_wishbone_bd_ram_n17805, p_wishbone_bd_ram_n17806,
         p_wishbone_bd_ram_n17807, p_wishbone_bd_ram_n17808,
         p_wishbone_bd_ram_n17809, p_wishbone_bd_ram_n17810,
         p_wishbone_bd_ram_n17811, p_wishbone_bd_ram_n17812,
         p_wishbone_bd_ram_n17813, p_wishbone_bd_ram_n17814,
         p_wishbone_bd_ram_n17815, p_wishbone_bd_ram_n17816,
         p_wishbone_bd_ram_n17817, p_wishbone_bd_ram_n17818,
         p_wishbone_bd_ram_n17819, p_wishbone_bd_ram_n17820,
         p_wishbone_bd_ram_n17821, p_wishbone_bd_ram_n17822,
         p_wishbone_bd_ram_n17823, p_wishbone_bd_ram_n17824,
         p_wishbone_bd_ram_n17825, p_wishbone_bd_ram_n17826,
         p_wishbone_bd_ram_n17827, p_wishbone_bd_ram_n17828,
         p_wishbone_bd_ram_n17829, p_wishbone_bd_ram_n17830,
         p_wishbone_bd_ram_n17831, p_wishbone_bd_ram_n17832,
         p_wishbone_bd_ram_n17833, p_wishbone_bd_ram_n17834,
         p_wishbone_bd_ram_n17835, p_wishbone_bd_ram_n17836,
         p_wishbone_bd_ram_n17837, p_wishbone_bd_ram_n17838,
         p_wishbone_bd_ram_n17839, p_wishbone_bd_ram_n17840,
         p_wishbone_bd_ram_n17841, p_wishbone_bd_ram_n17842,
         p_wishbone_bd_ram_n17843, p_wishbone_bd_ram_n17844,
         p_wishbone_bd_ram_n17845, p_wishbone_bd_ram_n17846,
         p_wishbone_bd_ram_n17847, p_wishbone_bd_ram_n17848,
         p_wishbone_bd_ram_n17849, p_wishbone_bd_ram_n17850,
         p_wishbone_bd_ram_n17851, p_wishbone_bd_ram_n17852,
         p_wishbone_bd_ram_n17853, p_wishbone_bd_ram_n17854,
         p_wishbone_bd_ram_n17855, p_wishbone_bd_ram_n17856,
         p_wishbone_bd_ram_n17857, p_wishbone_bd_ram_n17858,
         p_wishbone_bd_ram_n17859, p_wishbone_bd_ram_n17860,
         p_wishbone_bd_ram_n17861, p_wishbone_bd_ram_n17862,
         p_wishbone_bd_ram_n17863, p_wishbone_bd_ram_n17864,
         p_wishbone_bd_ram_n17865, p_wishbone_bd_ram_n17866,
         p_wishbone_bd_ram_n17867, p_wishbone_bd_ram_n17868,
         p_wishbone_bd_ram_n17869, p_wishbone_bd_ram_n17870,
         p_wishbone_bd_ram_n17871, p_wishbone_bd_ram_n17872,
         p_wishbone_bd_ram_n17873, p_wishbone_bd_ram_n17874,
         p_wishbone_bd_ram_n17875, p_wishbone_bd_ram_n17876,
         p_wishbone_bd_ram_n17877, p_wishbone_bd_ram_n17878,
         p_wishbone_bd_ram_n17879, p_wishbone_bd_ram_n17880,
         p_wishbone_bd_ram_n17881, p_wishbone_bd_ram_n17882,
         p_wishbone_bd_ram_n17883, p_wishbone_bd_ram_n17884,
         p_wishbone_bd_ram_n17885, p_wishbone_bd_ram_n17886,
         p_wishbone_bd_ram_n17887, p_wishbone_bd_ram_n17888,
         p_wishbone_bd_ram_n17889, p_wishbone_bd_ram_n17890,
         p_wishbone_bd_ram_n17891, p_wishbone_bd_ram_n17892,
         p_wishbone_bd_ram_n17893, p_wishbone_bd_ram_n17894,
         p_wishbone_bd_ram_n17895, p_wishbone_bd_ram_n17896,
         p_wishbone_bd_ram_n17897, p_wishbone_bd_ram_n17898,
         p_wishbone_bd_ram_n17899, p_wishbone_bd_ram_n17900,
         p_wishbone_bd_ram_n17901, p_wishbone_bd_ram_n17902,
         p_wishbone_bd_ram_n17903, p_wishbone_bd_ram_n17904,
         p_wishbone_bd_ram_n17905, p_wishbone_bd_ram_n17906,
         p_wishbone_bd_ram_n17907, p_wishbone_bd_ram_n17908,
         p_wishbone_bd_ram_n17909, p_wishbone_bd_ram_n17910,
         p_wishbone_bd_ram_n17911, p_wishbone_bd_ram_n17912,
         p_wishbone_bd_ram_n17913, p_wishbone_bd_ram_n17914,
         p_wishbone_bd_ram_n17915, p_wishbone_bd_ram_n17916,
         p_wishbone_bd_ram_n17917, p_wishbone_bd_ram_n17918,
         p_wishbone_bd_ram_n17919, p_wishbone_bd_ram_n17920,
         p_wishbone_bd_ram_n17921, p_wishbone_bd_ram_n17922,
         p_wishbone_bd_ram_n17923, p_wishbone_bd_ram_n17924,
         p_wishbone_bd_ram_n17925, p_wishbone_bd_ram_n17926,
         p_wishbone_bd_ram_n17927, p_wishbone_bd_ram_n17928,
         p_wishbone_bd_ram_n17929, p_wishbone_bd_ram_n17930,
         p_wishbone_bd_ram_n17931, p_wishbone_bd_ram_n17932,
         p_wishbone_bd_ram_n17933, p_wishbone_bd_ram_n17934,
         p_wishbone_bd_ram_n17935, p_wishbone_bd_ram_n17936,
         p_wishbone_bd_ram_n17937, p_wishbone_bd_ram_n17938,
         p_wishbone_bd_ram_n17939, p_wishbone_bd_ram_n17940,
         p_wishbone_bd_ram_n17941, p_wishbone_bd_ram_n17942,
         p_wishbone_bd_ram_n17943, p_wishbone_bd_ram_n17944,
         p_wishbone_bd_ram_n17945, p_wishbone_bd_ram_n17946,
         p_wishbone_bd_ram_n17947, p_wishbone_bd_ram_n17948,
         p_wishbone_bd_ram_n17949, p_wishbone_bd_ram_n17950,
         p_wishbone_bd_ram_n17951, p_wishbone_bd_ram_n17952,
         p_wishbone_bd_ram_n17953, p_wishbone_bd_ram_n17954,
         p_wishbone_bd_ram_n17955, p_wishbone_bd_ram_n17956,
         p_wishbone_bd_ram_n17957, p_wishbone_bd_ram_n17958,
         p_wishbone_bd_ram_n17959, p_wishbone_bd_ram_n17960,
         p_wishbone_bd_ram_n17961, p_wishbone_bd_ram_n17962,
         p_wishbone_bd_ram_n17963, p_wishbone_bd_ram_n17964,
         p_wishbone_bd_ram_n17965, p_wishbone_bd_ram_n17966,
         p_wishbone_bd_ram_n17967, p_wishbone_bd_ram_n17968,
         p_wishbone_bd_ram_n17969, p_wishbone_bd_ram_n17970,
         p_wishbone_bd_ram_n17971, p_wishbone_bd_ram_n17972,
         p_wishbone_bd_ram_n17973, p_wishbone_bd_ram_n17974,
         p_wishbone_bd_ram_n17975, p_wishbone_bd_ram_n17976,
         p_wishbone_bd_ram_n17977, p_wishbone_bd_ram_n17978,
         p_wishbone_bd_ram_n17979, p_wishbone_bd_ram_n17980,
         p_wishbone_bd_ram_n17981, p_wishbone_bd_ram_n17982,
         p_wishbone_bd_ram_n17983, p_wishbone_bd_ram_n17984,
         p_wishbone_bd_ram_n17985, p_wishbone_bd_ram_n17986,
         p_wishbone_bd_ram_n17987, p_wishbone_bd_ram_n17988,
         p_wishbone_bd_ram_n17989, p_wishbone_bd_ram_n17990,
         p_wishbone_bd_ram_n17991, p_wishbone_bd_ram_n17992,
         p_wishbone_bd_ram_n17993, p_wishbone_bd_ram_n17994,
         p_wishbone_bd_ram_n17995, p_wishbone_bd_ram_n17996,
         p_wishbone_bd_ram_n17997, p_wishbone_bd_ram_n17998,
         p_wishbone_bd_ram_n17999, p_wishbone_bd_ram_n18000,
         p_wishbone_bd_ram_n18001, p_wishbone_bd_ram_n18002,
         p_wishbone_bd_ram_n18003, p_wishbone_bd_ram_n18004,
         p_wishbone_bd_ram_n18005, p_wishbone_bd_ram_n18006,
         p_wishbone_bd_ram_n18007, p_wishbone_bd_ram_n18008,
         p_wishbone_bd_ram_n18009, p_wishbone_bd_ram_n18010,
         p_wishbone_bd_ram_n18011, p_wishbone_bd_ram_n18012,
         p_wishbone_bd_ram_n18013, p_wishbone_bd_ram_n18014,
         p_wishbone_bd_ram_n18015, p_wishbone_bd_ram_n18016,
         p_wishbone_bd_ram_n18017, p_wishbone_bd_ram_n18018,
         p_wishbone_bd_ram_n18019, p_wishbone_bd_ram_n18020,
         p_wishbone_bd_ram_n18021, p_wishbone_bd_ram_n18022,
         p_wishbone_bd_ram_n18023, p_wishbone_bd_ram_n18024,
         p_wishbone_bd_ram_n18025, p_wishbone_bd_ram_n18026,
         p_wishbone_bd_ram_n18027, p_wishbone_bd_ram_n18028,
         p_wishbone_bd_ram_n18029, p_wishbone_bd_ram_n18030,
         p_wishbone_bd_ram_n18031, p_wishbone_bd_ram_n18032,
         p_wishbone_bd_ram_n18033, p_wishbone_bd_ram_n18034,
         p_wishbone_bd_ram_n18035, p_wishbone_bd_ram_n18036,
         p_wishbone_bd_ram_n18037, p_wishbone_bd_ram_n18038,
         p_wishbone_bd_ram_n18039, p_wishbone_bd_ram_n18040,
         p_wishbone_bd_ram_n18041, p_wishbone_bd_ram_n18042,
         p_wishbone_bd_ram_n18043, p_wishbone_bd_ram_n18044,
         p_wishbone_bd_ram_n18045, p_wishbone_bd_ram_n18046,
         p_wishbone_bd_ram_n18047, p_wishbone_bd_ram_n18048,
         p_wishbone_bd_ram_n18049, p_wishbone_bd_ram_n18050,
         p_wishbone_bd_ram_n18051, p_wishbone_bd_ram_n18052,
         p_wishbone_bd_ram_n18053, p_wishbone_bd_ram_n18054,
         p_wishbone_bd_ram_n18055, p_wishbone_bd_ram_n18056,
         p_wishbone_bd_ram_n18057, p_wishbone_bd_ram_n18058,
         p_wishbone_bd_ram_n18059, p_wishbone_bd_ram_n18060,
         p_wishbone_bd_ram_n18061, p_wishbone_bd_ram_n18062,
         p_wishbone_bd_ram_n18063, p_wishbone_bd_ram_n18064,
         p_wishbone_bd_ram_n18065, p_wishbone_bd_ram_n18066,
         p_wishbone_bd_ram_n18067, p_wishbone_bd_ram_n18068,
         p_wishbone_bd_ram_n18069, p_wishbone_bd_ram_n18070,
         p_wishbone_bd_ram_n18071, p_wishbone_bd_ram_n18072,
         p_wishbone_bd_ram_n18073, p_wishbone_bd_ram_n18074,
         p_wishbone_bd_ram_n18075, p_wishbone_bd_ram_n18076,
         p_wishbone_bd_ram_n18077, p_wishbone_bd_ram_n18078,
         p_wishbone_bd_ram_n18079, p_wishbone_bd_ram_n18080,
         p_wishbone_bd_ram_n18081, p_wishbone_bd_ram_n18082,
         p_wishbone_bd_ram_n18083, p_wishbone_bd_ram_n18084,
         p_wishbone_bd_ram_n18085, p_wishbone_bd_ram_n18086,
         p_wishbone_bd_ram_n18087, p_wishbone_bd_ram_n18088,
         p_wishbone_bd_ram_n18089, p_wishbone_bd_ram_n18090,
         p_wishbone_bd_ram_n18091, p_wishbone_bd_ram_n18092,
         p_wishbone_bd_ram_n18093, p_wishbone_bd_ram_n18094,
         p_wishbone_bd_ram_n18095, p_wishbone_bd_ram_n18096,
         p_wishbone_bd_ram_n18097, p_wishbone_bd_ram_n18098,
         p_wishbone_bd_ram_n18099, p_wishbone_bd_ram_n18100,
         p_wishbone_bd_ram_n18101, p_wishbone_bd_ram_n18102,
         p_wishbone_bd_ram_n18103, p_wishbone_bd_ram_n18104,
         p_wishbone_bd_ram_n18105, p_wishbone_bd_ram_n18106,
         p_wishbone_bd_ram_n18107, p_wishbone_bd_ram_n18108,
         p_wishbone_bd_ram_n18109, p_wishbone_bd_ram_n18110,
         p_wishbone_bd_ram_n18111, p_wishbone_bd_ram_n18112,
         p_wishbone_bd_ram_n18113, p_wishbone_bd_ram_n18114,
         p_wishbone_bd_ram_n18115, p_wishbone_bd_ram_n18116,
         p_wishbone_bd_ram_n18117, p_wishbone_bd_ram_n18118,
         p_wishbone_bd_ram_n18119, p_wishbone_bd_ram_n18120,
         p_wishbone_bd_ram_n18121, p_wishbone_bd_ram_n18122,
         p_wishbone_bd_ram_n18123, p_wishbone_bd_ram_n18124,
         p_wishbone_bd_ram_n18125, p_wishbone_bd_ram_n18126,
         p_wishbone_bd_ram_n18127, p_wishbone_bd_ram_n18128,
         p_wishbone_bd_ram_n18129, p_wishbone_bd_ram_n18130,
         p_wishbone_bd_ram_n18131, p_wishbone_bd_ram_n18132,
         p_wishbone_bd_ram_n18133, p_wishbone_bd_ram_n18134,
         p_wishbone_bd_ram_n18135, p_wishbone_bd_ram_n18136,
         p_wishbone_bd_ram_n18137, p_wishbone_bd_ram_n18138,
         p_wishbone_bd_ram_n18139, p_wishbone_bd_ram_n18140,
         p_wishbone_bd_ram_n18141, p_wishbone_bd_ram_n18142,
         p_wishbone_bd_ram_n18143, p_wishbone_bd_ram_n18144,
         p_wishbone_bd_ram_n18145, p_wishbone_bd_ram_n18146,
         p_wishbone_bd_ram_n18147, p_wishbone_bd_ram_n18148,
         p_wishbone_bd_ram_n18149, p_wishbone_bd_ram_n18150,
         p_wishbone_bd_ram_n18151, p_wishbone_bd_ram_n18152,
         p_wishbone_bd_ram_n18153, p_wishbone_bd_ram_n18154,
         p_wishbone_bd_ram_n18155, p_wishbone_bd_ram_n18156,
         p_wishbone_bd_ram_n18157, p_wishbone_bd_ram_n18158,
         p_wishbone_bd_ram_n18159, p_wishbone_bd_ram_n18160,
         p_wishbone_bd_ram_n18161, p_wishbone_bd_ram_n18162,
         p_wishbone_bd_ram_n18163, p_wishbone_bd_ram_n18164,
         p_wishbone_bd_ram_n18165, p_wishbone_bd_ram_n18166,
         p_wishbone_bd_ram_n18167, p_wishbone_bd_ram_n18168,
         p_wishbone_bd_ram_n18169, p_wishbone_bd_ram_n18170,
         p_wishbone_bd_ram_n18171, p_wishbone_bd_ram_n18172,
         p_wishbone_bd_ram_n18173, p_wishbone_bd_ram_n18174,
         p_wishbone_bd_ram_n18175, p_wishbone_bd_ram_n18176,
         p_wishbone_bd_ram_n18177, p_wishbone_bd_ram_n18178,
         p_wishbone_bd_ram_n18179, p_wishbone_bd_ram_n18180,
         p_wishbone_bd_ram_n18181, p_wishbone_bd_ram_n18182,
         p_wishbone_bd_ram_n18183, p_wishbone_bd_ram_n18184,
         p_wishbone_bd_ram_n18185, p_wishbone_bd_ram_n18186,
         p_wishbone_bd_ram_n18187, p_wishbone_bd_ram_n18188,
         p_wishbone_bd_ram_n18189, p_wishbone_bd_ram_n18190,
         p_wishbone_bd_ram_n18191, p_wishbone_bd_ram_n18192,
         p_wishbone_bd_ram_n18193, p_wishbone_bd_ram_n18194,
         p_wishbone_bd_ram_n18195, p_wishbone_bd_ram_n18196,
         p_wishbone_bd_ram_n18197, p_wishbone_bd_ram_n18198,
         p_wishbone_bd_ram_n18199, p_wishbone_bd_ram_n18200,
         p_wishbone_bd_ram_n18201, p_wishbone_bd_ram_n18202,
         p_wishbone_bd_ram_n18203, p_wishbone_bd_ram_n18204,
         p_wishbone_bd_ram_n18205, p_wishbone_bd_ram_n18206,
         p_wishbone_bd_ram_n18207, p_wishbone_bd_ram_n18208,
         p_wishbone_bd_ram_n18209, p_wishbone_bd_ram_n18210,
         p_wishbone_bd_ram_n18211, p_wishbone_bd_ram_n18212,
         p_wishbone_bd_ram_n18213, p_wishbone_bd_ram_n18214,
         p_wishbone_bd_ram_n18215, p_wishbone_bd_ram_n18216,
         p_wishbone_bd_ram_n18217, p_wishbone_bd_ram_n18218,
         p_wishbone_bd_ram_n18219, p_wishbone_bd_ram_n18220,
         p_wishbone_bd_ram_n18221, p_wishbone_bd_ram_n18222,
         p_wishbone_bd_ram_n18223, p_wishbone_bd_ram_n18224,
         p_wishbone_bd_ram_n18225, p_wishbone_bd_ram_n18226,
         p_wishbone_bd_ram_n18227, p_wishbone_bd_ram_n18228,
         p_wishbone_bd_ram_n18229, p_wishbone_bd_ram_n18230,
         p_wishbone_bd_ram_n18231, p_wishbone_bd_ram_n18232,
         p_wishbone_bd_ram_n18233, p_wishbone_bd_ram_n18234,
         p_wishbone_bd_ram_n18235, p_wishbone_bd_ram_n18236,
         p_wishbone_bd_ram_n18237, p_wishbone_bd_ram_n18238,
         p_wishbone_bd_ram_n18239, p_wishbone_bd_ram_n18240,
         p_wishbone_bd_ram_n18241, p_wishbone_bd_ram_n18242,
         p_wishbone_bd_ram_n18243, p_wishbone_bd_ram_n18244,
         p_wishbone_bd_ram_n18245, p_wishbone_bd_ram_n18246,
         p_wishbone_bd_ram_n18247, p_wishbone_bd_ram_n18248,
         p_wishbone_bd_ram_n18249, p_wishbone_bd_ram_n18250,
         p_wishbone_bd_ram_n18251, p_wishbone_bd_ram_n18252,
         p_wishbone_bd_ram_n18253, p_wishbone_bd_ram_n18254,
         p_wishbone_bd_ram_n18255, p_wishbone_bd_ram_n18256,
         p_wishbone_bd_ram_n18257, p_wishbone_bd_ram_n18258,
         p_wishbone_bd_ram_n18259, p_wishbone_bd_ram_n18260,
         p_wishbone_bd_ram_n18261, p_wishbone_bd_ram_n18262,
         p_wishbone_bd_ram_n18263, p_wishbone_bd_ram_n18264,
         p_wishbone_bd_ram_n18265, p_wishbone_bd_ram_n18266,
         p_wishbone_bd_ram_n18267, p_wishbone_bd_ram_n18268,
         p_wishbone_bd_ram_n18269, p_wishbone_bd_ram_n18270,
         p_wishbone_bd_ram_n18271, p_wishbone_bd_ram_n18272,
         p_wishbone_bd_ram_n18273, p_wishbone_bd_ram_n18274,
         p_wishbone_bd_ram_n18275, p_wishbone_bd_ram_n18276,
         p_wishbone_bd_ram_n18277, p_wishbone_bd_ram_n18278,
         p_wishbone_bd_ram_n18279, p_wishbone_bd_ram_n18280,
         p_wishbone_bd_ram_n18281, p_wishbone_bd_ram_n18282,
         p_wishbone_bd_ram_n18283, p_wishbone_bd_ram_n18284,
         p_wishbone_bd_ram_n18285, p_wishbone_bd_ram_n18286,
         p_wishbone_bd_ram_n18287, p_wishbone_bd_ram_n18288,
         p_wishbone_bd_ram_n18289, p_wishbone_bd_ram_n18290,
         p_wishbone_bd_ram_n18291, p_wishbone_bd_ram_n18292,
         p_wishbone_bd_ram_n18293, p_wishbone_bd_ram_n18294,
         p_wishbone_bd_ram_n18295, p_wishbone_bd_ram_n18296,
         p_wishbone_bd_ram_n18297, p_wishbone_bd_ram_n18298,
         p_wishbone_bd_ram_n18299, p_wishbone_bd_ram_n18300,
         p_wishbone_bd_ram_n18301, p_wishbone_bd_ram_n18302,
         p_wishbone_bd_ram_n18303, p_wishbone_bd_ram_n18304,
         p_wishbone_bd_ram_n18305, p_wishbone_bd_ram_n18306,
         p_wishbone_bd_ram_n18307, p_wishbone_bd_ram_n18308,
         p_wishbone_bd_ram_n18309, p_wishbone_bd_ram_n18310,
         p_wishbone_bd_ram_n18311, p_wishbone_bd_ram_n18312,
         p_wishbone_bd_ram_n18313, p_wishbone_bd_ram_n18314,
         p_wishbone_bd_ram_n18315, p_wishbone_bd_ram_n18316,
         p_wishbone_bd_ram_n18317, p_wishbone_bd_ram_n18318,
         p_wishbone_bd_ram_n18319, p_wishbone_bd_ram_n18320,
         p_wishbone_bd_ram_n18321, p_wishbone_bd_ram_n18322,
         p_wishbone_bd_ram_n18323, p_wishbone_bd_ram_n18324,
         p_wishbone_bd_ram_n18325, p_wishbone_bd_ram_n18326,
         p_wishbone_bd_ram_n18327, p_wishbone_bd_ram_n18328,
         p_wishbone_bd_ram_n18329, p_wishbone_bd_ram_n18330,
         p_wishbone_bd_ram_n18331, p_wishbone_bd_ram_n18332,
         p_wishbone_bd_ram_n18333, p_wishbone_bd_ram_n18334,
         p_wishbone_bd_ram_n18335, p_wishbone_bd_ram_n18336,
         p_wishbone_bd_ram_n18337, p_wishbone_bd_ram_n18338,
         p_wishbone_bd_ram_n18339, p_wishbone_bd_ram_n18340,
         p_wishbone_bd_ram_n18341, p_wishbone_bd_ram_n18342,
         p_wishbone_bd_ram_n18343, p_wishbone_bd_ram_n18344,
         p_wishbone_bd_ram_n18345, p_wishbone_bd_ram_n18346,
         p_wishbone_bd_ram_n18347, p_wishbone_bd_ram_n18348,
         p_wishbone_bd_ram_n18349, p_wishbone_bd_ram_n18350,
         p_wishbone_bd_ram_n18351, p_wishbone_bd_ram_n18352,
         p_wishbone_bd_ram_n18353, p_wishbone_bd_ram_n18354,
         p_wishbone_bd_ram_n18355, p_wishbone_bd_ram_n18356,
         p_wishbone_bd_ram_n18357, p_wishbone_bd_ram_n18358,
         p_wishbone_bd_ram_n18359, p_wishbone_bd_ram_n18360,
         p_wishbone_bd_ram_n18361, p_wishbone_bd_ram_n18362,
         p_wishbone_bd_ram_n18363, p_wishbone_bd_ram_n18364,
         p_wishbone_bd_ram_n18365, p_wishbone_bd_ram_n18366,
         p_wishbone_bd_ram_n18367, p_wishbone_bd_ram_n18368,
         p_wishbone_bd_ram_n18369, p_wishbone_bd_ram_n18370,
         p_wishbone_bd_ram_n18371, p_wishbone_bd_ram_n18372,
         p_wishbone_bd_ram_n18373, p_wishbone_bd_ram_n18374,
         p_wishbone_bd_ram_n18375, p_wishbone_bd_ram_n18376,
         p_wishbone_bd_ram_n18377, p_wishbone_bd_ram_n18378,
         p_wishbone_bd_ram_n18379, p_wishbone_bd_ram_n18380,
         p_wishbone_bd_ram_n18381, p_wishbone_bd_ram_n18382,
         p_wishbone_bd_ram_n18383, p_wishbone_bd_ram_n18384,
         p_wishbone_bd_ram_n18385, p_wishbone_bd_ram_n18386,
         p_wishbone_bd_ram_n18387, p_wishbone_bd_ram_n18388,
         p_wishbone_bd_ram_n18389, p_wishbone_bd_ram_n18390,
         p_wishbone_bd_ram_n18391, p_wishbone_bd_ram_n18392,
         p_wishbone_bd_ram_n18393, p_wishbone_bd_ram_n18394,
         p_wishbone_bd_ram_n18395, p_wishbone_bd_ram_n18396,
         p_wishbone_bd_ram_n18397, p_wishbone_bd_ram_n18398,
         p_wishbone_bd_ram_n18399, p_wishbone_bd_ram_n18400,
         p_wishbone_bd_ram_n18401, p_wishbone_bd_ram_n18402,
         p_wishbone_bd_ram_n18403, p_wishbone_bd_ram_n18404,
         p_wishbone_bd_ram_n18405, p_wishbone_bd_ram_n18406,
         p_wishbone_bd_ram_n18407, p_wishbone_bd_ram_n18408,
         p_wishbone_bd_ram_n18409, p_wishbone_bd_ram_n18410,
         p_wishbone_bd_ram_n18411, p_wishbone_bd_ram_n18412,
         p_wishbone_bd_ram_n18413, p_wishbone_bd_ram_n18414,
         p_wishbone_bd_ram_n18415, p_wishbone_bd_ram_n18416,
         p_wishbone_bd_ram_n18417, p_wishbone_bd_ram_n18418,
         p_wishbone_bd_ram_n18419, p_wishbone_bd_ram_n18420,
         p_wishbone_bd_ram_n18421, p_wishbone_bd_ram_n18422,
         p_wishbone_bd_ram_n18423, p_wishbone_bd_ram_n18424,
         p_wishbone_bd_ram_n18425, p_wishbone_bd_ram_n18426,
         p_wishbone_bd_ram_n18427, p_wishbone_bd_ram_n18428,
         p_wishbone_bd_ram_n18429, p_wishbone_bd_ram_n18430,
         p_wishbone_bd_ram_n18431, p_wishbone_bd_ram_n18432,
         p_wishbone_bd_ram_n18433, p_wishbone_bd_ram_n18434,
         p_wishbone_bd_ram_n18435, p_wishbone_bd_ram_n18436,
         p_wishbone_bd_ram_n18437, p_wishbone_bd_ram_n18438,
         p_wishbone_bd_ram_n18439, p_wishbone_bd_ram_n18440,
         p_wishbone_bd_ram_n18441, p_wishbone_bd_ram_n18442,
         p_wishbone_bd_ram_n18443, p_wishbone_bd_ram_n18444,
         p_wishbone_bd_ram_n18445, p_wishbone_bd_ram_n18446,
         p_wishbone_bd_ram_n18447, p_wishbone_bd_ram_n18448,
         p_wishbone_bd_ram_n18449, p_wishbone_bd_ram_n18450,
         p_wishbone_bd_ram_n18451, p_wishbone_bd_ram_n18452,
         p_wishbone_bd_ram_n18453, p_wishbone_bd_ram_n18454,
         p_wishbone_bd_ram_n18455, p_wishbone_bd_ram_n18456,
         p_wishbone_bd_ram_n18457, p_wishbone_bd_ram_n18458,
         p_wishbone_bd_ram_n18459, p_wishbone_bd_ram_n18460,
         p_wishbone_bd_ram_n18461, p_wishbone_bd_ram_n18462,
         p_wishbone_bd_ram_n18463, p_wishbone_bd_ram_n18464,
         p_wishbone_bd_ram_n18465, p_wishbone_bd_ram_n18466,
         p_wishbone_bd_ram_n18467, p_wishbone_bd_ram_n18468,
         p_wishbone_bd_ram_n18469, p_wishbone_bd_ram_n18470,
         p_wishbone_bd_ram_n18471, p_wishbone_bd_ram_n18472,
         p_wishbone_bd_ram_n18473, p_wishbone_bd_ram_n18474,
         p_wishbone_bd_ram_n18475, p_wishbone_bd_ram_n18476,
         p_wishbone_bd_ram_n18477, p_wishbone_bd_ram_n18478,
         p_wishbone_bd_ram_n18479, p_wishbone_bd_ram_n18480,
         p_wishbone_bd_ram_n18481, p_wishbone_bd_ram_n18482,
         p_wishbone_bd_ram_n18483, p_wishbone_bd_ram_n18484,
         p_wishbone_bd_ram_n18485, p_wishbone_bd_ram_n18486,
         p_wishbone_bd_ram_n18487, p_wishbone_bd_ram_n18488,
         p_wishbone_bd_ram_n18489, p_wishbone_bd_ram_n18490,
         p_wishbone_bd_ram_n18491, p_wishbone_bd_ram_n18492,
         p_wishbone_bd_ram_n18493, p_wishbone_bd_ram_n18494,
         p_wishbone_bd_ram_n18495, p_wishbone_bd_ram_n18496,
         p_wishbone_bd_ram_n18497, p_wishbone_bd_ram_n18498,
         p_wishbone_bd_ram_n18499, p_wishbone_bd_ram_n18500,
         p_wishbone_bd_ram_n18501, p_wishbone_bd_ram_n18502,
         p_wishbone_bd_ram_n18503, p_wishbone_bd_ram_n18504,
         p_wishbone_bd_ram_n18505, p_wishbone_bd_ram_n18506,
         p_wishbone_bd_ram_n18507, p_wishbone_bd_ram_n18508,
         p_wishbone_bd_ram_n18509, p_wishbone_bd_ram_n18510,
         p_wishbone_bd_ram_n18511, p_wishbone_bd_ram_n18512,
         p_wishbone_bd_ram_n18513, p_wishbone_bd_ram_n18514,
         p_wishbone_bd_ram_n18515, p_wishbone_bd_ram_n18516,
         p_wishbone_bd_ram_n18517, p_wishbone_bd_ram_n18518,
         p_wishbone_bd_ram_n18519, p_wishbone_bd_ram_n18520,
         p_wishbone_bd_ram_n18521, p_wishbone_bd_ram_n18522,
         p_wishbone_bd_ram_n18523, p_wishbone_bd_ram_n18524,
         p_wishbone_bd_ram_n18525, p_wishbone_bd_ram_n18526,
         p_wishbone_bd_ram_n18527, p_wishbone_bd_ram_n18528,
         p_wishbone_bd_ram_n18529, p_wishbone_bd_ram_n18530,
         p_wishbone_bd_ram_n18531, p_wishbone_bd_ram_n18532,
         p_wishbone_bd_ram_n18533, p_wishbone_bd_ram_n18534,
         p_wishbone_bd_ram_n18535, p_wishbone_bd_ram_n18536,
         p_wishbone_bd_ram_n18537, p_wishbone_bd_ram_n18538,
         p_wishbone_bd_ram_n18539, p_wishbone_bd_ram_n18540,
         p_wishbone_bd_ram_n18541, p_wishbone_bd_ram_n18542,
         p_wishbone_bd_ram_n18543, p_wishbone_bd_ram_n18544,
         p_wishbone_bd_ram_n18545, p_wishbone_bd_ram_n18546,
         p_wishbone_bd_ram_n18547, p_wishbone_bd_ram_n18548,
         p_wishbone_bd_ram_n18549, p_wishbone_bd_ram_n18550,
         p_wishbone_bd_ram_n18551, p_wishbone_bd_ram_n18552,
         p_wishbone_bd_ram_n18553, p_wishbone_bd_ram_n18554,
         p_wishbone_bd_ram_n18555, p_wishbone_bd_ram_n18556,
         p_wishbone_bd_ram_n18557, p_wishbone_bd_ram_n18558,
         p_wishbone_bd_ram_n18559, p_wishbone_bd_ram_n18560,
         p_wishbone_bd_ram_n18561, p_wishbone_bd_ram_n18562,
         p_wishbone_bd_ram_n18563, p_wishbone_bd_ram_n18564,
         p_wishbone_bd_ram_n18565, p_wishbone_bd_ram_n18566,
         p_wishbone_bd_ram_n18567, p_wishbone_bd_ram_n18568,
         p_wishbone_bd_ram_n18569, p_wishbone_bd_ram_n18570,
         p_wishbone_bd_ram_n18571, p_wishbone_bd_ram_n18572,
         p_wishbone_bd_ram_n18573, p_wishbone_bd_ram_n18574,
         p_wishbone_bd_ram_n18575, p_wishbone_bd_ram_n18576,
         p_wishbone_bd_ram_n18577, p_wishbone_bd_ram_n18578,
         p_wishbone_bd_ram_n18579, p_wishbone_bd_ram_n18580,
         p_wishbone_bd_ram_n18581, p_wishbone_bd_ram_n18582,
         p_wishbone_bd_ram_n18583, p_wishbone_bd_ram_n18584,
         p_wishbone_bd_ram_n18585, p_wishbone_bd_ram_n18586,
         p_wishbone_bd_ram_n18587, p_wishbone_bd_ram_n18588,
         p_wishbone_bd_ram_n18589, p_wishbone_bd_ram_n18590,
         p_wishbone_bd_ram_n18591, p_wishbone_bd_ram_n18592,
         p_wishbone_bd_ram_n18593, p_wishbone_bd_ram_n18594,
         p_wishbone_bd_ram_n18595, p_wishbone_bd_ram_n18596,
         p_wishbone_bd_ram_n18597, p_wishbone_bd_ram_n18598,
         p_wishbone_bd_ram_n18599, p_wishbone_bd_ram_n18600,
         p_wishbone_bd_ram_n18601, p_wishbone_bd_ram_n18602,
         p_wishbone_bd_ram_n18603, p_wishbone_bd_ram_n18604,
         p_wishbone_bd_ram_n18605, p_wishbone_bd_ram_n18606,
         p_wishbone_bd_ram_n18607, p_wishbone_bd_ram_n18608,
         p_wishbone_bd_ram_n18609, p_wishbone_bd_ram_n18610,
         p_wishbone_bd_ram_n18611, p_wishbone_bd_ram_n18612,
         p_wishbone_bd_ram_n18613, p_wishbone_bd_ram_n18614,
         p_wishbone_bd_ram_n18615, p_wishbone_bd_ram_n18616,
         p_wishbone_bd_ram_n18617, p_wishbone_bd_ram_n18618,
         p_wishbone_bd_ram_n18619, p_wishbone_bd_ram_n18620,
         p_wishbone_bd_ram_n18621, p_wishbone_bd_ram_n18622,
         p_wishbone_bd_ram_n18623, p_wishbone_bd_ram_n18624,
         p_wishbone_bd_ram_n18625, p_wishbone_bd_ram_n18626,
         p_wishbone_bd_ram_n18627, p_wishbone_bd_ram_n18628,
         p_wishbone_bd_ram_n18629, p_wishbone_bd_ram_n18630,
         p_wishbone_bd_ram_n18631, p_wishbone_bd_ram_n18632,
         p_wishbone_bd_ram_n18633, p_wishbone_bd_ram_n18634,
         p_wishbone_bd_ram_n18635, p_wishbone_bd_ram_n18636,
         p_wishbone_bd_ram_n18637, p_wishbone_bd_ram_n18638,
         p_wishbone_bd_ram_n18639, p_wishbone_bd_ram_n18640,
         p_wishbone_bd_ram_n18641, p_wishbone_bd_ram_n18642,
         p_wishbone_bd_ram_n18643, p_wishbone_bd_ram_n18644,
         p_wishbone_bd_ram_n18645, p_wishbone_bd_ram_n18646,
         p_wishbone_bd_ram_n18647, p_wishbone_bd_ram_n18648,
         p_wishbone_bd_ram_n18649, p_wishbone_bd_ram_n18650,
         p_wishbone_bd_ram_n18651, p_wishbone_bd_ram_n18652,
         p_wishbone_bd_ram_n18653, p_wishbone_bd_ram_n18654,
         p_wishbone_bd_ram_n18655, p_wishbone_bd_ram_n18656,
         p_wishbone_bd_ram_n18657, p_wishbone_bd_ram_n18658,
         p_wishbone_bd_ram_n18659, p_wishbone_bd_ram_n18660,
         p_wishbone_bd_ram_n18661, p_wishbone_bd_ram_n18662,
         p_wishbone_bd_ram_n18663, p_wishbone_bd_ram_n18664,
         p_wishbone_bd_ram_n18665, p_wishbone_bd_ram_n18666,
         p_wishbone_bd_ram_n18667, p_wishbone_bd_ram_n18668,
         p_wishbone_bd_ram_n18669, p_wishbone_bd_ram_n18670,
         p_wishbone_bd_ram_n18671, p_wishbone_bd_ram_n18672,
         p_wishbone_bd_ram_n18673, p_wishbone_bd_ram_n18674,
         p_wishbone_bd_ram_n18675, p_wishbone_bd_ram_n18676,
         p_wishbone_bd_ram_n18677, p_wishbone_bd_ram_n18678,
         p_wishbone_bd_ram_n18679, p_wishbone_bd_ram_n18680,
         p_wishbone_bd_ram_n18681, p_wishbone_bd_ram_n18682,
         p_wishbone_bd_ram_n18683, p_wishbone_bd_ram_n18684,
         p_wishbone_bd_ram_n18685, p_wishbone_bd_ram_n18686,
         p_wishbone_bd_ram_n18687, p_wishbone_bd_ram_n18688,
         p_wishbone_bd_ram_n18689, p_wishbone_bd_ram_n18690,
         p_wishbone_bd_ram_n18691, p_wishbone_bd_ram_n18692,
         p_wishbone_bd_ram_n18693, p_wishbone_bd_ram_n18694,
         p_wishbone_bd_ram_n18695, p_wishbone_bd_ram_n18696,
         p_wishbone_bd_ram_n18697, p_wishbone_bd_ram_n18698,
         p_wishbone_bd_ram_n18699, p_wishbone_bd_ram_n18700,
         p_wishbone_bd_ram_n18701, p_wishbone_bd_ram_n18702,
         p_wishbone_bd_ram_n18703, p_wishbone_bd_ram_n18704,
         p_wishbone_bd_ram_n18705, p_wishbone_bd_ram_n18706,
         p_wishbone_bd_ram_n18707, p_wishbone_bd_ram_n18708,
         p_wishbone_bd_ram_n18709, p_wishbone_bd_ram_n18710,
         p_wishbone_bd_ram_n18711, p_wishbone_bd_ram_n18712,
         p_wishbone_bd_ram_n18713, p_wishbone_bd_ram_n18714,
         p_wishbone_bd_ram_n18715, p_wishbone_bd_ram_n18716,
         p_wishbone_bd_ram_n18717, p_wishbone_bd_ram_n18718,
         p_wishbone_bd_ram_n18719, p_wishbone_bd_ram_n18720,
         p_wishbone_bd_ram_n18721, p_wishbone_bd_ram_n18722,
         p_wishbone_bd_ram_n18723, p_wishbone_bd_ram_n18724,
         p_wishbone_bd_ram_n18725, p_wishbone_bd_ram_n18726,
         p_wishbone_bd_ram_n18727, p_wishbone_bd_ram_n18728,
         p_wishbone_bd_ram_n18729, p_wishbone_bd_ram_n18730,
         p_wishbone_bd_ram_n18731, p_wishbone_bd_ram_n18732,
         p_wishbone_bd_ram_n18733, p_wishbone_bd_ram_n18734,
         p_wishbone_bd_ram_n18735, p_wishbone_bd_ram_n18736,
         p_wishbone_bd_ram_n18737, p_wishbone_bd_ram_n18738,
         p_wishbone_bd_ram_n18739, p_wishbone_bd_ram_n18740,
         p_wishbone_bd_ram_n18741, p_wishbone_bd_ram_n18742,
         p_wishbone_bd_ram_n18743, p_wishbone_bd_ram_n18744,
         p_wishbone_bd_ram_n18745, p_wishbone_bd_ram_n18746,
         p_wishbone_bd_ram_n18747, p_wishbone_bd_ram_n18748,
         p_wishbone_bd_ram_n18749, p_wishbone_bd_ram_n18750,
         p_wishbone_bd_ram_n18751, p_wishbone_bd_ram_n18752,
         p_wishbone_bd_ram_n18753, p_wishbone_bd_ram_n18754,
         p_wishbone_bd_ram_n18755, p_wishbone_bd_ram_n18756,
         p_wishbone_bd_ram_n18757, p_wishbone_bd_ram_n18758,
         p_wishbone_bd_ram_n18759, p_wishbone_bd_ram_n18760,
         p_wishbone_bd_ram_n18761, p_wishbone_bd_ram_n18762,
         p_wishbone_bd_ram_n18763, p_wishbone_bd_ram_n18764,
         p_wishbone_bd_ram_n18765, p_wishbone_bd_ram_n18766,
         p_wishbone_bd_ram_n18767, p_wishbone_bd_ram_n18768,
         p_wishbone_bd_ram_n18769, p_wishbone_bd_ram_n18770,
         p_wishbone_bd_ram_n18771, p_wishbone_bd_ram_n18772,
         p_wishbone_bd_ram_n18773, p_wishbone_bd_ram_n18774,
         p_wishbone_bd_ram_n18775, p_wishbone_bd_ram_n18776,
         p_wishbone_bd_ram_n18777, p_wishbone_bd_ram_n18778,
         p_wishbone_bd_ram_n18779, p_wishbone_bd_ram_n18780,
         p_wishbone_bd_ram_n18781, p_wishbone_bd_ram_n18782,
         p_wishbone_bd_ram_n18783, p_wishbone_bd_ram_n18784,
         p_wishbone_bd_ram_n18785, p_wishbone_bd_ram_n18786,
         p_wishbone_bd_ram_n18787, p_wishbone_bd_ram_n18788,
         p_wishbone_bd_ram_n18789, p_wishbone_bd_ram_n18790,
         p_wishbone_bd_ram_n18791, p_wishbone_bd_ram_n18792,
         p_wishbone_bd_ram_n18793, p_wishbone_bd_ram_n18794,
         p_wishbone_bd_ram_n18795, p_wishbone_bd_ram_n18796,
         p_wishbone_bd_ram_n18797, p_wishbone_bd_ram_n18798,
         p_wishbone_bd_ram_n18799, p_wishbone_bd_ram_n18800,
         p_wishbone_bd_ram_n18801, p_wishbone_bd_ram_n18802,
         p_wishbone_bd_ram_n18803, p_wishbone_bd_ram_n18804,
         p_wishbone_bd_ram_n18805, p_wishbone_bd_ram_n18806,
         p_wishbone_bd_ram_n18807, p_wishbone_bd_ram_n18808,
         p_wishbone_bd_ram_n18809, p_wishbone_bd_ram_n18810,
         p_wishbone_bd_ram_n18811, p_wishbone_bd_ram_n18812,
         p_wishbone_bd_ram_n18813, p_wishbone_bd_ram_n18814,
         p_wishbone_bd_ram_n18815, p_wishbone_bd_ram_n18816,
         p_wishbone_bd_ram_n18817, p_wishbone_bd_ram_n18818,
         p_wishbone_bd_ram_n18819, p_wishbone_bd_ram_n18820,
         p_wishbone_bd_ram_n18821, p_wishbone_bd_ram_n18822,
         p_wishbone_bd_ram_n18823, p_wishbone_bd_ram_n18824,
         p_wishbone_bd_ram_n18825, p_wishbone_bd_ram_n18826,
         p_wishbone_bd_ram_n18827, p_wishbone_bd_ram_n18828,
         p_wishbone_bd_ram_n18829, p_wishbone_bd_ram_n18830,
         p_wishbone_bd_ram_n18831, p_wishbone_bd_ram_n18832,
         p_wishbone_bd_ram_n18833, p_wishbone_bd_ram_n18834,
         p_wishbone_bd_ram_n18835, p_wishbone_bd_ram_n18836,
         p_wishbone_bd_ram_n18837, p_wishbone_bd_ram_n18838,
         p_wishbone_bd_ram_n18839, p_wishbone_bd_ram_n18840,
         p_wishbone_bd_ram_n18841, p_wishbone_bd_ram_n18842,
         p_wishbone_bd_ram_n18843, p_wishbone_bd_ram_n18844,
         p_wishbone_bd_ram_n18845, p_wishbone_bd_ram_n18846,
         p_wishbone_bd_ram_n18847, p_wishbone_bd_ram_n18848,
         p_wishbone_bd_ram_n18849, p_wishbone_bd_ram_n18850,
         p_wishbone_bd_ram_n18851, p_wishbone_bd_ram_n18852,
         p_wishbone_bd_ram_n18853, p_wishbone_bd_ram_n18854,
         p_wishbone_bd_ram_n18855, p_wishbone_bd_ram_n18856,
         p_wishbone_bd_ram_n18857, p_wishbone_bd_ram_n18858,
         p_wishbone_bd_ram_n18859, p_wishbone_bd_ram_n18860,
         p_wishbone_bd_ram_n18861, p_wishbone_bd_ram_n18862,
         p_wishbone_bd_ram_n18863, p_wishbone_bd_ram_n18864,
         p_wishbone_bd_ram_n18865, p_wishbone_bd_ram_n18866,
         p_wishbone_bd_ram_n18867, p_wishbone_bd_ram_n18868,
         p_wishbone_bd_ram_n18869, p_wishbone_bd_ram_n18870,
         p_wishbone_bd_ram_n18871, p_wishbone_bd_ram_n18872,
         p_wishbone_bd_ram_n18873, p_wishbone_bd_ram_n18874,
         p_wishbone_bd_ram_n18875, p_wishbone_bd_ram_n18876,
         p_wishbone_bd_ram_n18877, p_wishbone_bd_ram_n18878,
         p_wishbone_bd_ram_n18879, p_wishbone_bd_ram_n18880,
         p_wishbone_bd_ram_n18881, p_wishbone_bd_ram_n18882,
         p_wishbone_bd_ram_n18883, p_wishbone_bd_ram_n18884,
         p_wishbone_bd_ram_n18885, p_wishbone_bd_ram_n18886,
         p_wishbone_bd_ram_n18887, p_wishbone_bd_ram_n18888,
         p_wishbone_bd_ram_n18889, p_wishbone_bd_ram_n18890,
         p_wishbone_bd_ram_n18891, p_wishbone_bd_ram_n18892,
         p_wishbone_bd_ram_n18893, p_wishbone_bd_ram_n18894,
         p_wishbone_bd_ram_n18895, p_wishbone_bd_ram_n18896,
         p_wishbone_bd_ram_n18897, p_wishbone_bd_ram_n18898,
         p_wishbone_bd_ram_n18899, p_wishbone_bd_ram_n18900,
         p_wishbone_bd_ram_n18901, p_wishbone_bd_ram_n18902,
         p_wishbone_bd_ram_n18903, p_wishbone_bd_ram_n18904,
         p_wishbone_bd_ram_n18905, p_wishbone_bd_ram_n18906,
         p_wishbone_bd_ram_n18907, p_wishbone_bd_ram_n18908,
         p_wishbone_bd_ram_n18909, p_wishbone_bd_ram_n18910,
         p_wishbone_bd_ram_n18911, p_wishbone_bd_ram_n18912,
         p_wishbone_bd_ram_n18913, p_wishbone_bd_ram_n18914,
         p_wishbone_bd_ram_n18915, p_wishbone_bd_ram_n18916,
         p_wishbone_bd_ram_n18917, p_wishbone_bd_ram_n18918,
         p_wishbone_bd_ram_n18919, p_wishbone_bd_ram_n18920,
         p_wishbone_bd_ram_n18921, p_wishbone_bd_ram_n18922,
         p_wishbone_bd_ram_n18923, p_wishbone_bd_ram_n18924,
         p_wishbone_bd_ram_n18925, p_wishbone_bd_ram_n18926,
         p_wishbone_bd_ram_n18927, p_wishbone_bd_ram_n18928,
         p_wishbone_bd_ram_n18929, p_wishbone_bd_ram_n18930,
         p_wishbone_bd_ram_n18931, p_wishbone_bd_ram_n18932,
         p_wishbone_bd_ram_n18933, p_wishbone_bd_ram_n18934,
         p_wishbone_bd_ram_n18935, p_wishbone_bd_ram_n18936,
         p_wishbone_bd_ram_n18937, p_wishbone_bd_ram_n18938,
         p_wishbone_bd_ram_n18939, p_wishbone_bd_ram_n18940,
         p_wishbone_bd_ram_n18941, p_wishbone_bd_ram_n18942,
         p_wishbone_bd_ram_n18943, p_wishbone_bd_ram_n18944,
         p_wishbone_bd_ram_n18945, p_wishbone_bd_ram_n18946,
         p_wishbone_bd_ram_n18947, p_wishbone_bd_ram_n18948,
         p_wishbone_bd_ram_n18949, p_wishbone_bd_ram_n18950,
         p_wishbone_bd_ram_n18951, p_wishbone_bd_ram_n18952,
         p_wishbone_bd_ram_n18953, p_wishbone_bd_ram_n18954,
         p_wishbone_bd_ram_n18955, p_wishbone_bd_ram_n18956,
         p_wishbone_bd_ram_n18957, p_wishbone_bd_ram_n18958,
         p_wishbone_bd_ram_n18959, p_wishbone_bd_ram_n18960,
         p_wishbone_bd_ram_n18961, p_wishbone_bd_ram_n18962,
         p_wishbone_bd_ram_n18963, p_wishbone_bd_ram_n18964,
         p_wishbone_bd_ram_n18965, p_wishbone_bd_ram_n18966,
         p_wishbone_bd_ram_n18967, p_wishbone_bd_ram_n18968,
         p_wishbone_bd_ram_n18969, p_wishbone_bd_ram_n18970,
         p_wishbone_bd_ram_n18971, p_wishbone_bd_ram_n18972,
         p_wishbone_bd_ram_n18973, p_wishbone_bd_ram_n18974,
         p_wishbone_bd_ram_n18975, p_wishbone_bd_ram_n18976,
         p_wishbone_bd_ram_n18977, p_wishbone_bd_ram_n18978,
         p_wishbone_bd_ram_n18979, p_wishbone_bd_ram_n18980,
         p_wishbone_bd_ram_n18981, p_wishbone_bd_ram_n18982,
         p_wishbone_bd_ram_n18983, p_wishbone_bd_ram_n18984,
         p_wishbone_bd_ram_n18985, p_wishbone_bd_ram_n18986,
         p_wishbone_bd_ram_n18987, p_wishbone_bd_ram_n18988,
         p_wishbone_bd_ram_n18989, p_wishbone_bd_ram_n18990,
         p_wishbone_bd_ram_n18991, p_wishbone_bd_ram_n18992,
         p_wishbone_bd_ram_n18993, p_wishbone_bd_ram_n18994,
         p_wishbone_bd_ram_n18995, p_wishbone_bd_ram_n18996,
         p_wishbone_bd_ram_n18997, p_wishbone_bd_ram_n18998,
         p_wishbone_bd_ram_n18999, p_wishbone_bd_ram_n19000,
         p_wishbone_bd_ram_n19001, p_wishbone_bd_ram_n19002,
         p_wishbone_bd_ram_n19003, p_wishbone_bd_ram_n19004,
         p_wishbone_bd_ram_n19005, p_wishbone_bd_ram_n19006,
         p_wishbone_bd_ram_n19007, p_wishbone_bd_ram_n19008,
         p_wishbone_bd_ram_n19009, p_wishbone_bd_ram_n19010,
         p_wishbone_bd_ram_n19011, p_wishbone_bd_ram_n19012,
         p_wishbone_bd_ram_n19013, p_wishbone_bd_ram_n19014,
         p_wishbone_bd_ram_n19015, p_wishbone_bd_ram_n19016,
         p_wishbone_bd_ram_n19017, p_wishbone_bd_ram_n19018,
         p_wishbone_bd_ram_n19019, p_wishbone_bd_ram_n19020,
         p_wishbone_bd_ram_n19021, p_wishbone_bd_ram_n19022,
         p_wishbone_bd_ram_n19023, p_wishbone_bd_ram_n19024,
         p_wishbone_bd_ram_n19025, p_wishbone_bd_ram_n19026,
         p_wishbone_bd_ram_n19027, p_wishbone_bd_ram_n19028,
         p_wishbone_bd_ram_n19029, p_wishbone_bd_ram_n19030,
         p_wishbone_bd_ram_n19031, p_wishbone_bd_ram_n19032,
         p_wishbone_bd_ram_n19033, p_wishbone_bd_ram_n19034,
         p_wishbone_bd_ram_n19035, p_wishbone_bd_ram_n19036,
         p_wishbone_bd_ram_n19037, p_wishbone_bd_ram_n19038,
         p_wishbone_bd_ram_n19039, p_wishbone_bd_ram_n19040,
         p_wishbone_bd_ram_n19041, p_wishbone_bd_ram_n19042,
         p_wishbone_bd_ram_n19043, p_wishbone_bd_ram_n19044,
         p_wishbone_bd_ram_n19045, p_wishbone_bd_ram_n19046,
         p_wishbone_bd_ram_n19047, p_wishbone_bd_ram_n19048,
         p_wishbone_bd_ram_n19049, p_wishbone_bd_ram_n19050,
         p_wishbone_bd_ram_n19051, p_wishbone_bd_ram_n19052,
         p_wishbone_bd_ram_n19053, p_wishbone_bd_ram_n19054,
         p_wishbone_bd_ram_n19055, p_wishbone_bd_ram_n19056,
         p_wishbone_bd_ram_n19057, p_wishbone_bd_ram_n19058,
         p_wishbone_bd_ram_n19059, p_wishbone_bd_ram_n19060,
         p_wishbone_bd_ram_n19061, p_wishbone_bd_ram_n19062,
         p_wishbone_bd_ram_n19063, p_wishbone_bd_ram_n19064,
         p_wishbone_bd_ram_n19065, p_wishbone_bd_ram_n19066,
         p_wishbone_bd_ram_n19067, p_wishbone_bd_ram_n19068,
         p_wishbone_bd_ram_n19069, p_wishbone_bd_ram_n19070,
         p_wishbone_bd_ram_n19071, p_wishbone_bd_ram_n19072,
         p_wishbone_bd_ram_n19073, p_wishbone_bd_ram_n19074,
         p_wishbone_bd_ram_n19075, p_wishbone_bd_ram_n19076,
         p_wishbone_bd_ram_n19077, p_wishbone_bd_ram_n19078,
         p_wishbone_bd_ram_n19079, p_wishbone_bd_ram_n19080,
         p_wishbone_bd_ram_n19081, p_wishbone_bd_ram_n19082,
         p_wishbone_bd_ram_n19083, p_wishbone_bd_ram_n19084,
         p_wishbone_bd_ram_n19085, p_wishbone_bd_ram_n19086,
         p_wishbone_bd_ram_n19087, p_wishbone_bd_ram_n19088,
         p_wishbone_bd_ram_n19089, p_wishbone_bd_ram_n19090,
         p_wishbone_bd_ram_n19091, p_wishbone_bd_ram_n19092,
         p_wishbone_bd_ram_n19093, p_wishbone_bd_ram_n19094,
         p_wishbone_bd_ram_n19095, p_wishbone_bd_ram_n19096,
         p_wishbone_bd_ram_n19097, p_wishbone_bd_ram_n19098,
         p_wishbone_bd_ram_n19099, p_wishbone_bd_ram_n19100,
         p_wishbone_bd_ram_n19101, p_wishbone_bd_ram_n19102,
         p_wishbone_bd_ram_n19103, p_wishbone_bd_ram_n19104,
         p_wishbone_bd_ram_n19105, p_wishbone_bd_ram_n19106,
         p_wishbone_bd_ram_n19107, p_wishbone_bd_ram_n19108,
         p_wishbone_bd_ram_n19109, p_wishbone_bd_ram_n19110,
         p_wishbone_bd_ram_n19111, p_wishbone_bd_ram_n19112,
         p_wishbone_bd_ram_n19113, p_wishbone_bd_ram_n19114,
         p_wishbone_bd_ram_n19115, p_wishbone_bd_ram_n19116,
         p_wishbone_bd_ram_n19117, p_wishbone_bd_ram_n19118,
         p_wishbone_bd_ram_n19119, p_wishbone_bd_ram_n19120,
         p_wishbone_bd_ram_n19121, p_wishbone_bd_ram_n19122,
         p_wishbone_bd_ram_n19123, p_wishbone_bd_ram_n19124,
         p_wishbone_bd_ram_n19125, p_wishbone_bd_ram_n19126,
         p_wishbone_bd_ram_n19127, p_wishbone_bd_ram_n19128,
         p_wishbone_bd_ram_n19129, p_wishbone_bd_ram_n19130,
         p_wishbone_bd_ram_n19131, p_wishbone_bd_ram_n19132,
         p_wishbone_bd_ram_n19133, p_wishbone_bd_ram_n19134,
         p_wishbone_bd_ram_n19135, p_wishbone_bd_ram_n19136,
         p_wishbone_bd_ram_n19137, p_wishbone_bd_ram_n19138,
         p_wishbone_bd_ram_n19139, p_wishbone_bd_ram_n19140,
         p_wishbone_bd_ram_n19141, p_wishbone_bd_ram_n19142,
         p_wishbone_bd_ram_n19143, p_wishbone_bd_ram_n19144,
         p_wishbone_bd_ram_n19145, p_wishbone_bd_ram_n19146,
         p_wishbone_bd_ram_n19147, p_wishbone_bd_ram_n19148,
         p_wishbone_bd_ram_n19149, p_wishbone_bd_ram_n19150,
         p_wishbone_bd_ram_n19151, p_wishbone_bd_ram_n19152,
         p_wishbone_bd_ram_n19153, p_wishbone_bd_ram_n19154,
         p_wishbone_bd_ram_n19155, p_wishbone_bd_ram_n19156,
         p_wishbone_bd_ram_n19157, p_wishbone_bd_ram_n19158,
         p_wishbone_bd_ram_n19159, p_wishbone_bd_ram_n19160,
         p_wishbone_bd_ram_n19161, p_wishbone_bd_ram_n19162,
         p_wishbone_bd_ram_n19163, p_wishbone_bd_ram_n19164,
         p_wishbone_bd_ram_n19165, p_wishbone_bd_ram_n19166,
         p_wishbone_bd_ram_n19167, p_wishbone_bd_ram_n19168,
         p_wishbone_bd_ram_n19169, p_wishbone_bd_ram_n19170,
         p_wishbone_bd_ram_n19171, p_wishbone_bd_ram_n19172,
         p_wishbone_bd_ram_n19173, p_wishbone_bd_ram_n19174,
         p_wishbone_bd_ram_n19175, p_wishbone_bd_ram_n19176,
         p_wishbone_bd_ram_n19177, p_wishbone_bd_ram_n19178,
         p_wishbone_bd_ram_n19179, p_wishbone_bd_ram_n19180,
         p_wishbone_bd_ram_n19181, p_wishbone_bd_ram_n19182,
         p_wishbone_bd_ram_n19183, p_wishbone_bd_ram_n19184,
         p_wishbone_bd_ram_n19185, p_wishbone_bd_ram_n19186,
         p_wishbone_bd_ram_n19187, p_wishbone_bd_ram_n19188,
         p_wishbone_bd_ram_n19189, p_wishbone_bd_ram_n19190,
         p_wishbone_bd_ram_n19191, p_wishbone_bd_ram_n19192,
         p_wishbone_bd_ram_n19193, p_wishbone_bd_ram_n19194,
         p_wishbone_bd_ram_n19195, p_wishbone_bd_ram_n19196,
         p_wishbone_bd_ram_n19197, p_wishbone_bd_ram_n19198,
         p_wishbone_bd_ram_n19199, p_wishbone_bd_ram_n19200,
         p_wishbone_bd_ram_n19201, p_wishbone_bd_ram_n19202,
         p_wishbone_bd_ram_n19203, p_wishbone_bd_ram_n19204,
         p_wishbone_bd_ram_n19205, p_wishbone_bd_ram_n19206,
         p_wishbone_bd_ram_n19207, p_wishbone_bd_ram_n19208,
         p_wishbone_bd_ram_n19209, p_wishbone_bd_ram_n19210,
         p_wishbone_bd_ram_n19211, p_wishbone_bd_ram_n19212,
         p_wishbone_bd_ram_n19213, p_wishbone_bd_ram_n19214,
         p_wishbone_bd_ram_n19215, p_wishbone_bd_ram_n19216,
         p_wishbone_bd_ram_n19217, p_wishbone_bd_ram_n19218,
         p_wishbone_bd_ram_n19219, p_wishbone_bd_ram_n19220,
         p_wishbone_bd_ram_n19221, p_wishbone_bd_ram_n19222,
         p_wishbone_bd_ram_n19223, p_wishbone_bd_ram_n19224,
         p_wishbone_bd_ram_n19225, p_wishbone_bd_ram_n19226,
         p_wishbone_bd_ram_n19227, p_wishbone_bd_ram_n19228,
         p_wishbone_bd_ram_n19229, p_wishbone_bd_ram_n19230,
         p_wishbone_bd_ram_n19231, p_wishbone_bd_ram_n19232,
         p_wishbone_bd_ram_n19233, p_wishbone_bd_ram_n19234,
         p_wishbone_bd_ram_n19235, p_wishbone_bd_ram_n19236,
         p_wishbone_bd_ram_n19237, p_wishbone_bd_ram_n19238,
         p_wishbone_bd_ram_n19239, p_wishbone_bd_ram_n19240,
         p_wishbone_bd_ram_n19241, p_wishbone_bd_ram_n19242,
         p_wishbone_bd_ram_n19243, p_wishbone_bd_ram_n19244,
         p_wishbone_bd_ram_n19245, p_wishbone_bd_ram_n19246,
         p_wishbone_bd_ram_n19247, p_wishbone_bd_ram_n19248,
         p_wishbone_bd_ram_n19249, p_wishbone_bd_ram_n19250,
         p_wishbone_bd_ram_n19251, p_wishbone_bd_ram_n19252,
         p_wishbone_bd_ram_n19253, p_wishbone_bd_ram_n19254,
         p_wishbone_bd_ram_n19255, p_wishbone_bd_ram_n19256,
         p_wishbone_bd_ram_n19257, p_wishbone_bd_ram_n19258,
         p_wishbone_bd_ram_n19259, p_wishbone_bd_ram_n19260,
         p_wishbone_bd_ram_n19261, p_wishbone_bd_ram_n19262,
         p_wishbone_bd_ram_n19263, p_wishbone_bd_ram_n19264,
         p_wishbone_bd_ram_n19265, p_wishbone_bd_ram_n19266,
         p_wishbone_bd_ram_n19267, p_wishbone_bd_ram_n19268,
         p_wishbone_bd_ram_n19269, p_wishbone_bd_ram_n19270,
         p_wishbone_bd_ram_n19271, p_wishbone_bd_ram_n19272,
         p_wishbone_bd_ram_n19273, p_wishbone_bd_ram_n19274,
         p_wishbone_bd_ram_n19275, p_wishbone_bd_ram_n19276,
         p_wishbone_bd_ram_n19277, p_wishbone_bd_ram_n19278,
         p_wishbone_bd_ram_n19279, p_wishbone_bd_ram_n19280,
         p_wishbone_bd_ram_n19281, p_wishbone_bd_ram_n19282,
         p_wishbone_bd_ram_n19283, p_wishbone_bd_ram_n19284,
         p_wishbone_bd_ram_n19285, p_wishbone_bd_ram_n19286,
         p_wishbone_bd_ram_n19287, p_wishbone_bd_ram_n19288,
         p_wishbone_bd_ram_n19289, p_wishbone_bd_ram_n19290,
         p_wishbone_bd_ram_n19291, p_wishbone_bd_ram_n19292,
         p_wishbone_bd_ram_n19293, p_wishbone_bd_ram_n19294,
         p_wishbone_bd_ram_n19295, p_wishbone_bd_ram_n19296,
         p_wishbone_bd_ram_n19297, p_wishbone_bd_ram_n19298,
         p_wishbone_bd_ram_n19299, p_wishbone_bd_ram_n19300,
         p_wishbone_bd_ram_n19301, p_wishbone_bd_ram_n19302,
         p_wishbone_bd_ram_n19303, p_wishbone_bd_ram_n19304,
         p_wishbone_bd_ram_n19305, p_wishbone_bd_ram_n19306,
         p_wishbone_bd_ram_n19307, p_wishbone_bd_ram_n19308,
         p_wishbone_bd_ram_n19309, p_wishbone_bd_ram_n19310,
         p_wishbone_bd_ram_n19311, p_wishbone_bd_ram_n19312,
         p_wishbone_bd_ram_n19313, p_wishbone_bd_ram_n19314,
         p_wishbone_bd_ram_n19315, p_wishbone_bd_ram_n19316,
         p_wishbone_bd_ram_n19317, p_wishbone_bd_ram_n19318,
         p_wishbone_bd_ram_n19319, p_wishbone_bd_ram_n19320,
         p_wishbone_bd_ram_n19321, p_wishbone_bd_ram_n19322,
         p_wishbone_bd_ram_n19323, p_wishbone_bd_ram_n19324,
         p_wishbone_bd_ram_n19325, p_wishbone_bd_ram_n19326,
         p_wishbone_bd_ram_n19327, p_wishbone_bd_ram_n19328,
         p_wishbone_bd_ram_n19329, p_wishbone_bd_ram_n19330,
         p_wishbone_bd_ram_n19331, p_wishbone_bd_ram_n19332,
         p_wishbone_bd_ram_n19333, p_wishbone_bd_ram_n19334,
         p_wishbone_bd_ram_n19335, p_wishbone_bd_ram_n19336,
         p_wishbone_bd_ram_n19337, p_wishbone_bd_ram_n19338,
         p_wishbone_bd_ram_n19339, p_wishbone_bd_ram_n19340,
         p_wishbone_bd_ram_n19341, p_wishbone_bd_ram_n19342,
         p_wishbone_bd_ram_n19343, p_wishbone_bd_ram_n19344,
         p_wishbone_bd_ram_n19345, p_wishbone_bd_ram_n19346,
         p_wishbone_bd_ram_n19347, p_wishbone_bd_ram_n19348,
         p_wishbone_bd_ram_n19349, p_wishbone_bd_ram_n19350,
         p_wishbone_bd_ram_n19351, p_wishbone_bd_ram_n19352,
         p_wishbone_bd_ram_n19353, p_wishbone_bd_ram_n19354,
         p_wishbone_bd_ram_n19355, p_wishbone_bd_ram_n19356,
         p_wishbone_bd_ram_n19357, p_wishbone_bd_ram_n19358,
         p_wishbone_bd_ram_n19359, p_wishbone_bd_ram_n19360,
         p_wishbone_bd_ram_n19361, p_wishbone_bd_ram_n19362,
         p_wishbone_bd_ram_n19363, p_wishbone_bd_ram_n19364,
         p_wishbone_bd_ram_n19365, p_wishbone_bd_ram_n19366,
         p_wishbone_bd_ram_n19367, p_wishbone_bd_ram_n19368,
         p_wishbone_bd_ram_n19369, p_wishbone_bd_ram_n19370,
         p_wishbone_bd_ram_n19371, p_wishbone_bd_ram_n19372,
         p_wishbone_bd_ram_n19373, p_wishbone_bd_ram_n19374,
         p_wishbone_bd_ram_n19375, p_wishbone_bd_ram_n19376,
         p_wishbone_bd_ram_n19377, p_wishbone_bd_ram_n19378,
         p_wishbone_bd_ram_n19379, p_wishbone_bd_ram_n19380,
         p_wishbone_bd_ram_n19381, p_wishbone_bd_ram_n19382,
         p_wishbone_bd_ram_n19383, p_wishbone_bd_ram_n19384,
         p_wishbone_bd_ram_n19385, p_wishbone_bd_ram_n19386,
         p_wishbone_bd_ram_n19387, p_wishbone_bd_ram_n19388,
         p_wishbone_bd_ram_n19389, p_wishbone_bd_ram_n19390,
         p_wishbone_bd_ram_n19391, p_wishbone_bd_ram_n19392,
         p_wishbone_bd_ram_n19393, p_wishbone_bd_ram_n19394,
         p_wishbone_bd_ram_n19395, p_wishbone_bd_ram_n19396,
         p_wishbone_bd_ram_n19397, p_wishbone_bd_ram_n19398,
         p_wishbone_bd_ram_n19399, p_wishbone_bd_ram_n19400,
         p_wishbone_bd_ram_n19401, p_wishbone_bd_ram_n19402,
         p_wishbone_bd_ram_n19403, p_wishbone_bd_ram_n19404,
         p_wishbone_bd_ram_n19405, p_wishbone_bd_ram_n19406,
         p_wishbone_bd_ram_n19407, p_wishbone_bd_ram_n19408,
         p_wishbone_bd_ram_n19409, p_wishbone_bd_ram_n19410,
         p_wishbone_bd_ram_n19411, p_wishbone_bd_ram_n19412,
         p_wishbone_bd_ram_n19413, p_wishbone_bd_ram_n19414,
         p_wishbone_bd_ram_n19415, p_wishbone_bd_ram_n19416,
         p_wishbone_bd_ram_n19417, p_wishbone_bd_ram_n19418,
         p_wishbone_bd_ram_n19419, p_wishbone_bd_ram_n19420,
         p_wishbone_bd_ram_n19421, p_wishbone_bd_ram_n19422,
         p_wishbone_bd_ram_n19423, p_wishbone_bd_ram_n19424,
         p_wishbone_bd_ram_n19425, p_wishbone_bd_ram_n19426,
         p_wishbone_bd_ram_n19427, p_wishbone_bd_ram_n19428,
         p_wishbone_bd_ram_n19429, p_wishbone_bd_ram_n19430,
         p_wishbone_bd_ram_n19431, p_wishbone_bd_ram_n19432,
         p_wishbone_bd_ram_n19433, p_wishbone_bd_ram_n19434,
         p_wishbone_bd_ram_n19435, p_wishbone_bd_ram_n19436,
         p_wishbone_bd_ram_n19437, p_wishbone_bd_ram_n19438,
         p_wishbone_bd_ram_n19439, p_wishbone_bd_ram_n19440,
         p_wishbone_bd_ram_n19441, p_wishbone_bd_ram_n19442,
         p_wishbone_bd_ram_n19443, p_wishbone_bd_ram_n19444,
         p_wishbone_bd_ram_n19445, p_wishbone_bd_ram_n19446,
         p_wishbone_bd_ram_n19447, p_wishbone_bd_ram_n19448,
         p_wishbone_bd_ram_n19449, p_wishbone_bd_ram_n19450,
         p_wishbone_bd_ram_n19451, p_wishbone_bd_ram_n19452,
         p_wishbone_bd_ram_n19453, p_wishbone_bd_ram_n19454,
         p_wishbone_bd_ram_n19455, p_wishbone_bd_ram_n19456,
         p_wishbone_bd_ram_n19457, p_wishbone_bd_ram_n19458,
         p_wishbone_bd_ram_n19459, p_wishbone_bd_ram_n19460,
         p_wishbone_bd_ram_n19461, p_wishbone_bd_ram_n19462,
         p_wishbone_bd_ram_n19463, p_wishbone_bd_ram_n19464,
         p_wishbone_bd_ram_n19465, p_wishbone_bd_ram_n19466,
         p_wishbone_bd_ram_n19467, p_wishbone_bd_ram_n19468,
         p_wishbone_bd_ram_n19469, p_wishbone_bd_ram_n19470,
         p_wishbone_bd_ram_n19471, p_wishbone_bd_ram_n19472,
         p_wishbone_bd_ram_n19473, p_wishbone_bd_ram_n19474,
         p_wishbone_bd_ram_n19475, p_wishbone_bd_ram_n19476,
         p_wishbone_bd_ram_n19477, p_wishbone_bd_ram_n19478,
         p_wishbone_bd_ram_n19479, p_wishbone_bd_ram_n19480,
         p_wishbone_bd_ram_n19481, p_wishbone_bd_ram_n19482,
         p_wishbone_bd_ram_n19483, p_wishbone_bd_ram_n19484,
         p_wishbone_bd_ram_n19485, p_wishbone_bd_ram_n19486,
         p_wishbone_bd_ram_n19487, p_wishbone_bd_ram_n19488,
         p_wishbone_bd_ram_n19489, p_wishbone_bd_ram_n19490,
         p_wishbone_bd_ram_n19491, p_wishbone_bd_ram_n19492,
         p_wishbone_bd_ram_n19493, p_wishbone_bd_ram_n19494,
         p_wishbone_bd_ram_n19495, p_wishbone_bd_ram_n19496,
         p_wishbone_bd_ram_n19497, p_wishbone_bd_ram_n19498,
         p_wishbone_bd_ram_n19499, p_wishbone_bd_ram_n19500,
         p_wishbone_bd_ram_n19501, p_wishbone_bd_ram_n19502,
         p_wishbone_bd_ram_n19503, p_wishbone_bd_ram_n19504,
         p_wishbone_bd_ram_n19505, p_wishbone_bd_ram_n19506,
         p_wishbone_bd_ram_n19507, p_wishbone_bd_ram_n19508,
         p_wishbone_bd_ram_n19509, p_wishbone_bd_ram_n19510,
         p_wishbone_bd_ram_n19511, p_wishbone_bd_ram_n19512,
         p_wishbone_bd_ram_n19513, p_wishbone_bd_ram_n19514,
         p_wishbone_bd_ram_n19515, p_wishbone_bd_ram_n19516,
         p_wishbone_bd_ram_n19517, p_wishbone_bd_ram_n19518,
         p_wishbone_bd_ram_n19519, p_wishbone_bd_ram_n19520,
         p_wishbone_bd_ram_n19521, p_wishbone_bd_ram_n19522,
         p_wishbone_bd_ram_n19523, p_wishbone_bd_ram_n19524,
         p_wishbone_bd_ram_n19525, p_wishbone_bd_ram_n19526,
         p_wishbone_bd_ram_n19527, p_wishbone_bd_ram_n19528,
         p_wishbone_bd_ram_n19529, p_wishbone_bd_ram_n19530,
         p_wishbone_bd_ram_n19531, p_wishbone_bd_ram_n19532,
         p_wishbone_bd_ram_n19533, p_wishbone_bd_ram_n19534,
         p_wishbone_bd_ram_n19535, p_wishbone_bd_ram_n19536,
         p_wishbone_bd_ram_n19537, p_wishbone_bd_ram_n19538,
         p_wishbone_bd_ram_n19539, p_wishbone_bd_ram_n19540,
         p_wishbone_bd_ram_n19541, p_wishbone_bd_ram_n19542,
         p_wishbone_bd_ram_n19543, p_wishbone_bd_ram_n19544,
         p_wishbone_bd_ram_n19545, p_wishbone_bd_ram_n19546,
         p_wishbone_bd_ram_n19547, p_wishbone_bd_ram_n19548,
         p_wishbone_bd_ram_n19549, p_wishbone_bd_ram_n19550,
         p_wishbone_bd_ram_n19551, p_wishbone_bd_ram_n19552,
         p_wishbone_bd_ram_n19553, p_wishbone_bd_ram_n19554,
         p_wishbone_bd_ram_n19555, p_wishbone_bd_ram_n19556,
         p_wishbone_bd_ram_n19557, p_wishbone_bd_ram_n19558,
         p_wishbone_bd_ram_n19559, p_wishbone_bd_ram_n19560,
         p_wishbone_bd_ram_n19561, p_wishbone_bd_ram_n19562,
         p_wishbone_bd_ram_n19563, p_wishbone_bd_ram_n19564,
         p_wishbone_bd_ram_n19565, p_wishbone_bd_ram_n19566,
         p_wishbone_bd_ram_n19567, p_wishbone_bd_ram_n19568,
         p_wishbone_bd_ram_n19569, p_wishbone_bd_ram_n19570,
         p_wishbone_bd_ram_n19571, p_wishbone_bd_ram_n19572,
         p_wishbone_bd_ram_n19573, p_wishbone_bd_ram_n19574,
         p_wishbone_bd_ram_n19575, p_wishbone_bd_ram_n19576,
         p_wishbone_bd_ram_n19577, p_wishbone_bd_ram_n19578,
         p_wishbone_bd_ram_n19579, p_wishbone_bd_ram_n19580,
         p_wishbone_bd_ram_n19581, p_wishbone_bd_ram_n19582,
         p_wishbone_bd_ram_n19583, p_wishbone_bd_ram_n19584,
         p_wishbone_bd_ram_n19585, p_wishbone_bd_ram_n19586,
         p_wishbone_bd_ram_n19587, p_wishbone_bd_ram_n19588,
         p_wishbone_bd_ram_n19589, p_wishbone_bd_ram_n19590,
         p_wishbone_bd_ram_n19591, p_wishbone_bd_ram_n19592,
         p_wishbone_bd_ram_n19593, p_wishbone_bd_ram_n19594,
         p_wishbone_bd_ram_n19595, p_wishbone_bd_ram_n19596,
         p_wishbone_bd_ram_n19597, p_wishbone_bd_ram_n19598,
         p_wishbone_bd_ram_n19599, p_wishbone_bd_ram_n19600,
         p_wishbone_bd_ram_n19601, p_wishbone_bd_ram_n19602,
         p_wishbone_bd_ram_n19603, p_wishbone_bd_ram_n19604,
         p_wishbone_bd_ram_n19605, p_wishbone_bd_ram_n19606,
         p_wishbone_bd_ram_n19607, p_wishbone_bd_ram_n19608,
         p_wishbone_bd_ram_n19609, p_wishbone_bd_ram_n19610,
         p_wishbone_bd_ram_n19611, p_wishbone_bd_ram_n19612,
         p_wishbone_bd_ram_n19613, p_wishbone_bd_ram_n19614,
         p_wishbone_bd_ram_n19615, p_wishbone_bd_ram_n19616,
         p_wishbone_bd_ram_n19617, p_wishbone_bd_ram_n19618,
         p_wishbone_bd_ram_n19619, p_wishbone_bd_ram_n19620,
         p_wishbone_bd_ram_n19621, p_wishbone_bd_ram_n19622,
         p_wishbone_bd_ram_n19623, p_wishbone_bd_ram_n19624,
         p_wishbone_bd_ram_n19625, p_wishbone_bd_ram_n19626,
         p_wishbone_bd_ram_n19627, p_wishbone_bd_ram_n19628,
         p_wishbone_bd_ram_n19629, p_wishbone_bd_ram_n19630,
         p_wishbone_bd_ram_n19631, p_wishbone_bd_ram_n19632,
         p_wishbone_bd_ram_n19633, p_wishbone_bd_ram_n19634,
         p_wishbone_bd_ram_n19635, p_wishbone_bd_ram_n19636,
         p_wishbone_bd_ram_n19637, p_wishbone_bd_ram_n19638,
         p_wishbone_bd_ram_n19639, p_wishbone_bd_ram_n19640,
         p_wishbone_bd_ram_n19641, p_wishbone_bd_ram_n19642,
         p_wishbone_bd_ram_n19643, p_wishbone_bd_ram_n19644,
         p_wishbone_bd_ram_n19645, p_wishbone_bd_ram_n19646,
         p_wishbone_bd_ram_n19647, p_wishbone_bd_ram_n19648,
         p_wishbone_bd_ram_n19649, p_wishbone_bd_ram_n19650,
         p_wishbone_bd_ram_n19651, p_wishbone_bd_ram_n19652,
         p_wishbone_bd_ram_n19653, p_wishbone_bd_ram_n19654,
         p_wishbone_bd_ram_n19655, p_wishbone_bd_ram_n19656,
         p_wishbone_bd_ram_n19657, p_wishbone_bd_ram_n19658,
         p_wishbone_bd_ram_n19659, p_wishbone_bd_ram_n19660,
         p_wishbone_bd_ram_n19661, p_wishbone_bd_ram_n19662,
         p_wishbone_bd_ram_n19663, p_wishbone_bd_ram_n19664,
         p_wishbone_bd_ram_n19665, p_wishbone_bd_ram_n19666,
         p_wishbone_bd_ram_n19667, p_wishbone_bd_ram_n19668,
         p_wishbone_bd_ram_n19669, p_wishbone_bd_ram_n19670,
         p_wishbone_bd_ram_n19671, p_wishbone_bd_ram_n19672,
         p_wishbone_bd_ram_n19673, p_wishbone_bd_ram_n19674,
         p_wishbone_bd_ram_n19675, p_wishbone_bd_ram_n19676,
         p_wishbone_bd_ram_n19677, p_wishbone_bd_ram_n19678,
         p_wishbone_bd_ram_n19679, p_wishbone_bd_ram_n19680,
         p_wishbone_bd_ram_n19681, p_wishbone_bd_ram_n19682,
         p_wishbone_bd_ram_n19683, p_wishbone_bd_ram_n19684,
         p_wishbone_bd_ram_n19685, p_wishbone_bd_ram_n19686,
         p_wishbone_bd_ram_n19687, p_wishbone_bd_ram_n19688,
         p_wishbone_bd_ram_n19689, p_wishbone_bd_ram_n19690,
         p_wishbone_bd_ram_n19691, p_wishbone_bd_ram_n19692,
         p_wishbone_bd_ram_n19693, p_wishbone_bd_ram_n19694,
         p_wishbone_bd_ram_n19695, p_wishbone_bd_ram_n19696,
         p_wishbone_bd_ram_n19697, p_wishbone_bd_ram_n19698,
         p_wishbone_bd_ram_n19699, p_wishbone_bd_ram_n19700,
         p_wishbone_bd_ram_n19701, p_wishbone_bd_ram_n19702,
         p_wishbone_bd_ram_n19703, p_wishbone_bd_ram_n19704,
         p_wishbone_bd_ram_n19705, p_wishbone_bd_ram_n19706,
         p_wishbone_bd_ram_n19707, p_wishbone_bd_ram_n19708,
         p_wishbone_bd_ram_n19709, p_wishbone_bd_ram_n19710,
         p_wishbone_bd_ram_n19711, p_wishbone_bd_ram_n19712,
         p_wishbone_bd_ram_n19713, p_wishbone_bd_ram_n19714,
         p_wishbone_bd_ram_n19715, p_wishbone_bd_ram_n19716,
         p_wishbone_bd_ram_n19717, p_wishbone_bd_ram_n19718,
         p_wishbone_bd_ram_n19719, p_wishbone_bd_ram_n19720,
         p_wishbone_bd_ram_n19721, p_wishbone_bd_ram_n19722,
         p_wishbone_bd_ram_n19723, p_wishbone_bd_ram_n19724,
         p_wishbone_bd_ram_n19725, p_wishbone_bd_ram_n19726,
         p_wishbone_bd_ram_n19727, p_wishbone_bd_ram_n19728,
         p_wishbone_bd_ram_n19729, p_wishbone_bd_ram_n19730,
         p_wishbone_bd_ram_n19731, p_wishbone_bd_ram_n19732,
         p_wishbone_bd_ram_n19733, p_wishbone_bd_ram_n19734,
         p_wishbone_bd_ram_n19735, p_wishbone_bd_ram_n19736,
         p_wishbone_bd_ram_n19737, p_wishbone_bd_ram_n19738,
         p_wishbone_bd_ram_n19739, p_wishbone_bd_ram_n19740,
         p_wishbone_bd_ram_n19741, p_wishbone_bd_ram_n19742,
         p_wishbone_bd_ram_n19743, p_wishbone_bd_ram_n19744,
         p_wishbone_bd_ram_n19745, p_wishbone_bd_ram_n19746,
         p_wishbone_bd_ram_n19747, p_wishbone_bd_ram_n19748,
         p_wishbone_bd_ram_n19749, p_wishbone_bd_ram_n19750,
         p_wishbone_bd_ram_n19751, p_wishbone_bd_ram_n19752,
         p_wishbone_bd_ram_n19753, p_wishbone_bd_ram_n19754,
         p_wishbone_bd_ram_n19755, p_wishbone_bd_ram_n19756,
         p_wishbone_bd_ram_n19757, p_wishbone_bd_ram_n19758,
         p_wishbone_bd_ram_n19759, p_wishbone_bd_ram_n19760,
         p_wishbone_bd_ram_n19761, p_wishbone_bd_ram_n19762,
         p_wishbone_bd_ram_n19763, p_wishbone_bd_ram_n19764,
         p_wishbone_bd_ram_n19765, p_wishbone_bd_ram_n19766,
         p_wishbone_bd_ram_n19767, p_wishbone_bd_ram_n19768,
         p_wishbone_bd_ram_n19769, p_wishbone_bd_ram_n19770,
         p_wishbone_bd_ram_n19771, p_wishbone_bd_ram_n19772,
         p_wishbone_bd_ram_n19773, p_wishbone_bd_ram_n19774,
         p_wishbone_bd_ram_n19775, p_wishbone_bd_ram_n19776,
         p_wishbone_bd_ram_n19777, p_wishbone_bd_ram_n19778,
         p_wishbone_bd_ram_n19779, p_wishbone_bd_ram_n19780,
         p_wishbone_bd_ram_n19781, p_wishbone_bd_ram_n19782,
         p_wishbone_bd_ram_n19783, p_wishbone_bd_ram_n19784,
         p_wishbone_bd_ram_n19785, p_wishbone_bd_ram_n19786,
         p_wishbone_bd_ram_n19787, p_wishbone_bd_ram_n19788,
         p_wishbone_bd_ram_n19789, p_wishbone_bd_ram_n19790,
         p_wishbone_bd_ram_n19791, p_wishbone_bd_ram_n19792,
         p_wishbone_bd_ram_n19793, p_wishbone_bd_ram_n19794,
         p_wishbone_bd_ram_n19795, p_wishbone_bd_ram_n19796,
         p_wishbone_bd_ram_n19797, p_wishbone_bd_ram_n19798,
         p_wishbone_bd_ram_n19799, p_wishbone_bd_ram_n19800,
         p_wishbone_bd_ram_n19801, p_wishbone_bd_ram_n19802,
         p_wishbone_bd_ram_n19803, p_wishbone_bd_ram_n19804,
         p_wishbone_bd_ram_n19805, p_wishbone_bd_ram_n19806,
         p_wishbone_bd_ram_n19807, p_wishbone_bd_ram_n19808,
         p_wishbone_bd_ram_n19809, p_wishbone_bd_ram_n19810,
         p_wishbone_bd_ram_n19811, p_wishbone_bd_ram_n19812,
         p_wishbone_bd_ram_n19813, p_wishbone_bd_ram_n19814,
         p_wishbone_bd_ram_n19815, p_wishbone_bd_ram_n19816,
         p_wishbone_bd_ram_n19817, p_wishbone_bd_ram_n19818,
         p_wishbone_bd_ram_n19819, p_wishbone_bd_ram_n19820,
         p_wishbone_bd_ram_n19821, p_wishbone_bd_ram_n19822,
         p_wishbone_bd_ram_n19823, p_wishbone_bd_ram_n19824,
         p_wishbone_bd_ram_n19825, p_wishbone_bd_ram_n19826,
         p_wishbone_bd_ram_n19827, p_wishbone_bd_ram_n19828,
         p_wishbone_bd_ram_n19829, p_wishbone_bd_ram_n19830,
         p_wishbone_bd_ram_n19831, p_wishbone_bd_ram_n19832,
         p_wishbone_bd_ram_n19833, p_wishbone_bd_ram_n19834,
         p_wishbone_bd_ram_n19835, p_wishbone_bd_ram_n19836,
         p_wishbone_bd_ram_n19837, p_wishbone_bd_ram_n19838,
         p_wishbone_bd_ram_n19839, p_wishbone_bd_ram_n19840,
         p_wishbone_bd_ram_n19841, p_wishbone_bd_ram_n19842,
         p_wishbone_bd_ram_n19843, p_wishbone_bd_ram_n19844,
         p_wishbone_bd_ram_n19845, p_wishbone_bd_ram_n19846,
         p_wishbone_bd_ram_n19847, p_wishbone_bd_ram_n19848,
         p_wishbone_bd_ram_n19849, p_wishbone_bd_ram_n19850,
         p_wishbone_bd_ram_n19851, p_wishbone_bd_ram_n19852,
         p_wishbone_bd_ram_n19853, p_wishbone_bd_ram_n19854,
         p_wishbone_bd_ram_n19855, p_wishbone_bd_ram_n19856,
         p_wishbone_bd_ram_n19857, p_wishbone_bd_ram_n19858,
         p_wishbone_bd_ram_n19859, p_wishbone_bd_ram_n19860,
         p_wishbone_bd_ram_n19861, p_wishbone_bd_ram_n19862,
         p_wishbone_bd_ram_n19863, p_wishbone_bd_ram_n19864,
         p_wishbone_bd_ram_n19865, p_wishbone_bd_ram_n19866,
         p_wishbone_bd_ram_n19867, p_wishbone_bd_ram_n19868,
         p_wishbone_bd_ram_n19869, p_wishbone_bd_ram_n19870,
         p_wishbone_bd_ram_n19871, p_wishbone_bd_ram_n19872,
         p_wishbone_bd_ram_n19873, p_wishbone_bd_ram_n19874,
         p_wishbone_bd_ram_n19875, p_wishbone_bd_ram_n19876,
         p_wishbone_bd_ram_n19877, p_wishbone_bd_ram_n19878,
         p_wishbone_bd_ram_n19879, p_wishbone_bd_ram_n19880,
         p_wishbone_bd_ram_n19881, p_wishbone_bd_ram_n19882,
         p_wishbone_bd_ram_n19883, p_wishbone_bd_ram_n19884,
         p_wishbone_bd_ram_n19885, p_wishbone_bd_ram_n19886,
         p_wishbone_bd_ram_n19887, p_wishbone_bd_ram_n19888,
         p_wishbone_bd_ram_n19889, p_wishbone_bd_ram_n19890,
         p_wishbone_bd_ram_n19891, p_wishbone_bd_ram_n19892,
         p_wishbone_bd_ram_n19893, p_wishbone_bd_ram_n19894,
         p_wishbone_bd_ram_n19895, p_wishbone_bd_ram_n19896,
         p_wishbone_bd_ram_n19897, p_wishbone_bd_ram_n19898,
         p_wishbone_bd_ram_n19899, p_wishbone_bd_ram_n19900,
         p_wishbone_bd_ram_n19901, p_wishbone_bd_ram_n19902,
         p_wishbone_bd_ram_n19903, p_wishbone_bd_ram_n19904,
         p_wishbone_bd_ram_n19905, p_wishbone_bd_ram_n19906,
         p_wishbone_bd_ram_n19907, p_wishbone_bd_ram_n19908,
         p_wishbone_bd_ram_n19909, p_wishbone_bd_ram_n19910,
         p_wishbone_bd_ram_n19911, p_wishbone_bd_ram_n19912,
         p_wishbone_bd_ram_n19913, p_wishbone_bd_ram_n19914,
         p_wishbone_bd_ram_n19915, p_wishbone_bd_ram_n19916,
         p_wishbone_bd_ram_n19917, p_wishbone_bd_ram_n19918,
         p_wishbone_bd_ram_n19919, p_wishbone_bd_ram_n19920,
         p_wishbone_bd_ram_n19921, p_wishbone_bd_ram_n19922,
         p_wishbone_bd_ram_n19923, p_wishbone_bd_ram_n19924,
         p_wishbone_bd_ram_n19925, p_wishbone_bd_ram_n19926,
         p_wishbone_bd_ram_n19927, p_wishbone_bd_ram_n19928,
         p_wishbone_bd_ram_n19929, p_wishbone_bd_ram_n19930,
         p_wishbone_bd_ram_n19931, p_wishbone_bd_ram_n19932,
         p_wishbone_bd_ram_n19933, p_wishbone_bd_ram_n19934,
         p_wishbone_bd_ram_n19935, p_wishbone_bd_ram_n19936,
         p_wishbone_bd_ram_n19937, p_wishbone_bd_ram_n19938,
         p_wishbone_bd_ram_n19939, p_wishbone_bd_ram_n19940,
         p_wishbone_bd_ram_n19941, p_wishbone_bd_ram_n19942,
         p_wishbone_bd_ram_n19943, p_wishbone_bd_ram_n19944,
         p_wishbone_bd_ram_n19945, p_wishbone_bd_ram_n19946,
         p_wishbone_bd_ram_n19947, p_wishbone_bd_ram_n19948,
         p_wishbone_bd_ram_n19949, p_wishbone_bd_ram_n19950,
         p_wishbone_bd_ram_n19951, p_wishbone_bd_ram_n19952,
         p_wishbone_bd_ram_n19953, p_wishbone_bd_ram_n19954,
         p_wishbone_bd_ram_n19955, p_wishbone_bd_ram_n19956,
         p_wishbone_bd_ram_n19957, p_wishbone_bd_ram_n19958,
         p_wishbone_bd_ram_n19959, p_wishbone_bd_ram_n19960,
         p_wishbone_bd_ram_n19961, p_wishbone_bd_ram_n19962,
         p_wishbone_bd_ram_n19963, p_wishbone_bd_ram_n19964,
         p_wishbone_bd_ram_n19965, p_wishbone_bd_ram_n19966,
         p_wishbone_bd_ram_n19967, p_wishbone_bd_ram_n19968,
         p_wishbone_bd_ram_n19969, p_wishbone_bd_ram_n19970,
         p_wishbone_bd_ram_n19971, p_wishbone_bd_ram_n19972,
         p_wishbone_bd_ram_n19973, p_wishbone_bd_ram_n19974,
         p_wishbone_bd_ram_n19975, p_wishbone_bd_ram_n19976,
         p_wishbone_bd_ram_n19977, p_wishbone_bd_ram_n19978,
         p_wishbone_bd_ram_n19979, p_wishbone_bd_ram_n19980,
         p_wishbone_bd_ram_n19981, p_wishbone_bd_ram_n19982,
         p_wishbone_bd_ram_n19983, p_wishbone_bd_ram_n19984,
         p_wishbone_bd_ram_n19985, p_wishbone_bd_ram_n19986,
         p_wishbone_bd_ram_n19987, p_wishbone_bd_ram_n19988,
         p_wishbone_bd_ram_n19989, p_wishbone_bd_ram_n19990,
         p_wishbone_bd_ram_n19991, p_wishbone_bd_ram_n19992,
         p_wishbone_bd_ram_n19993, p_wishbone_bd_ram_n19994,
         p_wishbone_bd_ram_n19995, p_wishbone_bd_ram_n19996,
         p_wishbone_bd_ram_n19997, p_wishbone_bd_ram_n19998,
         p_wishbone_bd_ram_n19999, p_wishbone_bd_ram_n20000,
         p_wishbone_bd_ram_n20001, p_wishbone_bd_ram_n20002,
         p_wishbone_bd_ram_n20003, p_wishbone_bd_ram_n20004,
         p_wishbone_bd_ram_n20005, p_wishbone_bd_ram_n20006,
         p_wishbone_bd_ram_n20007, p_wishbone_bd_ram_n20008,
         p_wishbone_bd_ram_n20009, p_wishbone_bd_ram_n20010,
         p_wishbone_bd_ram_n20011, p_wishbone_bd_ram_n20012,
         p_wishbone_bd_ram_n20013, p_wishbone_bd_ram_n20014,
         p_wishbone_bd_ram_n20015, p_wishbone_bd_ram_n20016,
         p_wishbone_bd_ram_n20017, p_wishbone_bd_ram_n20018,
         p_wishbone_bd_ram_n20019, p_wishbone_bd_ram_n20020,
         p_wishbone_bd_ram_n20021, p_wishbone_bd_ram_n20022,
         p_wishbone_bd_ram_n20023, p_wishbone_bd_ram_n20024,
         p_wishbone_bd_ram_n20025, p_wishbone_bd_ram_n20026,
         p_wishbone_bd_ram_n20027, p_wishbone_bd_ram_n20028,
         p_wishbone_bd_ram_n20029, p_wishbone_bd_ram_n20030,
         p_wishbone_bd_ram_n20031, p_wishbone_bd_ram_n20032,
         p_wishbone_bd_ram_n20033, p_wishbone_bd_ram_n20034,
         p_wishbone_bd_ram_n20035, p_wishbone_bd_ram_n20036,
         p_wishbone_bd_ram_n20037, p_wishbone_bd_ram_n20038,
         p_wishbone_bd_ram_n20039, p_wishbone_bd_ram_n20040,
         p_wishbone_bd_ram_n20041, p_wishbone_bd_ram_n20042,
         p_wishbone_bd_ram_n20043, p_wishbone_bd_ram_n20044,
         p_wishbone_bd_ram_n20045, p_wishbone_bd_ram_n20046,
         p_wishbone_bd_ram_n20047, p_wishbone_bd_ram_n20048,
         p_wishbone_bd_ram_n20049, p_wishbone_bd_ram_n20050,
         p_wishbone_bd_ram_n20051, p_wishbone_bd_ram_n20052,
         p_wishbone_bd_ram_n20053, p_wishbone_bd_ram_n20054,
         p_wishbone_bd_ram_n20055, p_wishbone_bd_ram_n20056,
         p_wishbone_bd_ram_n20057, p_wishbone_bd_ram_n20058,
         p_wishbone_bd_ram_n20059, p_wishbone_bd_ram_n20060,
         p_wishbone_bd_ram_n20061, p_wishbone_bd_ram_n20062,
         p_wishbone_bd_ram_n20063, p_wishbone_bd_ram_n20064,
         p_wishbone_bd_ram_n20065, p_wishbone_bd_ram_n20066,
         p_wishbone_bd_ram_n20067, p_wishbone_bd_ram_n20068,
         p_wishbone_bd_ram_n20069, p_wishbone_bd_ram_n20070,
         p_wishbone_bd_ram_n20071, p_wishbone_bd_ram_n20072,
         p_wishbone_bd_ram_n20073, p_wishbone_bd_ram_n20074,
         p_wishbone_bd_ram_n20075, p_wishbone_bd_ram_n20076,
         p_wishbone_bd_ram_n20077, p_wishbone_bd_ram_n20078,
         p_wishbone_bd_ram_n20079, p_wishbone_bd_ram_n20080,
         p_wishbone_bd_ram_n20081, p_wishbone_bd_ram_n20082,
         p_wishbone_bd_ram_n20083, p_wishbone_bd_ram_n20084,
         p_wishbone_bd_ram_n20085, p_wishbone_bd_ram_n20086,
         p_wishbone_bd_ram_n20087, p_wishbone_bd_ram_n20088,
         p_wishbone_bd_ram_n20089, p_wishbone_bd_ram_n20090,
         p_wishbone_bd_ram_n20091, p_wishbone_bd_ram_n20092,
         p_wishbone_bd_ram_n20093, p_wishbone_bd_ram_n20094,
         p_wishbone_bd_ram_n20095, p_wishbone_bd_ram_n20096,
         p_wishbone_bd_ram_n20097, p_wishbone_bd_ram_n20098,
         p_wishbone_bd_ram_n20099, p_wishbone_bd_ram_n20100,
         p_wishbone_bd_ram_n20101, p_wishbone_bd_ram_n20102,
         p_wishbone_bd_ram_n20103, p_wishbone_bd_ram_n20104,
         p_wishbone_bd_ram_n20105, p_wishbone_bd_ram_n20106,
         p_wishbone_bd_ram_n20107, p_wishbone_bd_ram_n20108,
         p_wishbone_bd_ram_n20109, p_wishbone_bd_ram_n20110,
         p_wishbone_bd_ram_n20111, p_wishbone_bd_ram_n20112,
         p_wishbone_bd_ram_n20113, p_wishbone_bd_ram_n20114,
         p_wishbone_bd_ram_n20115, p_wishbone_bd_ram_n20116,
         p_wishbone_bd_ram_n20117, p_wishbone_bd_ram_n20118,
         p_wishbone_bd_ram_n20119, p_wishbone_bd_ram_n20120,
         p_wishbone_bd_ram_n20121, p_wishbone_bd_ram_n20122,
         p_wishbone_bd_ram_n20123, p_wishbone_bd_ram_n20124,
         p_wishbone_bd_ram_n20125, p_wishbone_bd_ram_n20126,
         p_wishbone_bd_ram_n20127, p_wishbone_bd_ram_n20128,
         p_wishbone_bd_ram_n20129, p_wishbone_bd_ram_n20130,
         p_wishbone_bd_ram_n20131, p_wishbone_bd_ram_n20132,
         p_wishbone_bd_ram_n20133, p_wishbone_bd_ram_n20134,
         p_wishbone_bd_ram_n20135, p_wishbone_bd_ram_n20136,
         p_wishbone_bd_ram_n20137, p_wishbone_bd_ram_n20138,
         p_wishbone_bd_ram_n20139, p_wishbone_bd_ram_n20140,
         p_wishbone_bd_ram_n20141, p_wishbone_bd_ram_n20142,
         p_wishbone_bd_ram_n20143, p_wishbone_bd_ram_n20144,
         p_wishbone_bd_ram_n20145, p_wishbone_bd_ram_n20146,
         p_wishbone_bd_ram_n20147, p_wishbone_bd_ram_n20148,
         p_wishbone_bd_ram_n20149, p_wishbone_bd_ram_n20150,
         p_wishbone_bd_ram_n20151, p_wishbone_bd_ram_n20152,
         p_wishbone_bd_ram_n20153, p_wishbone_bd_ram_n20154,
         p_wishbone_bd_ram_n20155, p_wishbone_bd_ram_n20156,
         p_wishbone_bd_ram_n20157, p_wishbone_bd_ram_n20158,
         p_wishbone_bd_ram_n20159, p_wishbone_bd_ram_n20160,
         p_wishbone_bd_ram_n20161, p_wishbone_bd_ram_n20162,
         p_wishbone_bd_ram_n20163, p_wishbone_bd_ram_n20164,
         p_wishbone_bd_ram_n20165, p_wishbone_bd_ram_n20166,
         p_wishbone_bd_ram_n20167, p_wishbone_bd_ram_n20168,
         p_wishbone_bd_ram_n20169, p_wishbone_bd_ram_n20170,
         p_wishbone_bd_ram_n20171, p_wishbone_bd_ram_n20172,
         p_wishbone_bd_ram_n20173, p_wishbone_bd_ram_n20174,
         p_wishbone_bd_ram_n20175, p_wishbone_bd_ram_n20176,
         p_wishbone_bd_ram_n20177, p_wishbone_bd_ram_n20178,
         p_wishbone_bd_ram_n20179, p_wishbone_bd_ram_n20180,
         p_wishbone_bd_ram_n20181, p_wishbone_bd_ram_n20182,
         p_wishbone_bd_ram_n20183, p_wishbone_bd_ram_n20184,
         p_wishbone_bd_ram_n20185, p_wishbone_bd_ram_n20186,
         p_wishbone_bd_ram_n20187, p_wishbone_bd_ram_n20188,
         p_wishbone_bd_ram_n20189, p_wishbone_bd_ram_n20190,
         p_wishbone_bd_ram_n20191, p_wishbone_bd_ram_n20192,
         p_wishbone_bd_ram_n20193, p_wishbone_bd_ram_n20194,
         p_wishbone_bd_ram_n20195, p_wishbone_bd_ram_n20196,
         p_wishbone_bd_ram_n20197, p_wishbone_bd_ram_n20198,
         p_wishbone_bd_ram_n20199, p_wishbone_bd_ram_n20200,
         p_wishbone_bd_ram_n20201, p_wishbone_bd_ram_n20202,
         p_wishbone_bd_ram_n20203, p_wishbone_bd_ram_n20204,
         p_wishbone_bd_ram_n20205, p_wishbone_bd_ram_n20206,
         p_wishbone_bd_ram_n20207, p_wishbone_bd_ram_n20208,
         p_wishbone_bd_ram_n20209, p_wishbone_bd_ram_n20210,
         p_wishbone_bd_ram_n20211, p_wishbone_bd_ram_n20212,
         p_wishbone_bd_ram_n20213, p_wishbone_bd_ram_n20214,
         p_wishbone_bd_ram_n20215, p_wishbone_bd_ram_n20216,
         p_wishbone_bd_ram_n20217, p_wishbone_bd_ram_n20218,
         p_wishbone_bd_ram_n20219, p_wishbone_bd_ram_n20220,
         p_wishbone_bd_ram_n20221, p_wishbone_bd_ram_n20222,
         p_wishbone_bd_ram_n20223, p_wishbone_bd_ram_n20224,
         p_wishbone_bd_ram_n20225, p_wishbone_bd_ram_n20226,
         p_wishbone_bd_ram_n20227, p_wishbone_bd_ram_n20228,
         p_wishbone_bd_ram_n20229, p_wishbone_bd_ram_n20230,
         p_wishbone_bd_ram_n20231, p_wishbone_bd_ram_n20232,
         p_wishbone_bd_ram_n20233, p_wishbone_bd_ram_n20234,
         p_wishbone_bd_ram_n20235, p_wishbone_bd_ram_n20236,
         p_wishbone_bd_ram_n20237, p_wishbone_bd_ram_n20238,
         p_wishbone_bd_ram_n20239, p_wishbone_bd_ram_n20240,
         p_wishbone_bd_ram_n20241, p_wishbone_bd_ram_n20242,
         p_wishbone_bd_ram_n20243, p_wishbone_bd_ram_n20244,
         p_wishbone_bd_ram_n20245, p_wishbone_bd_ram_n20246,
         p_wishbone_bd_ram_n20247, p_wishbone_bd_ram_n20248,
         p_wishbone_bd_ram_n20249, p_wishbone_bd_ram_n20250,
         p_wishbone_bd_ram_n20251, p_wishbone_bd_ram_n20252,
         p_wishbone_bd_ram_n20253, p_wishbone_bd_ram_n20254,
         p_wishbone_bd_ram_n20255, p_wishbone_bd_ram_n20256,
         p_wishbone_bd_ram_n20257, p_wishbone_bd_ram_n20258,
         p_wishbone_bd_ram_n20259, p_wishbone_bd_ram_n20260,
         p_wishbone_bd_ram_n20261, p_wishbone_bd_ram_n20262,
         p_wishbone_bd_ram_n20263, p_wishbone_bd_ram_n20264,
         p_wishbone_bd_ram_n20265, p_wishbone_bd_ram_n20266,
         p_wishbone_bd_ram_n20267, p_wishbone_bd_ram_n20268,
         p_wishbone_bd_ram_n20269, p_wishbone_bd_ram_n20270,
         p_wishbone_bd_ram_n20271, p_wishbone_bd_ram_n20272,
         p_wishbone_bd_ram_n20273, p_wishbone_bd_ram_n20274,
         p_wishbone_bd_ram_n20275, p_wishbone_bd_ram_n20276,
         p_wishbone_bd_ram_n20277, p_wishbone_bd_ram_n20278,
         p_wishbone_bd_ram_n20279, p_wishbone_bd_ram_n20280,
         p_wishbone_bd_ram_n20281, p_wishbone_bd_ram_n20282,
         p_wishbone_bd_ram_n20283, p_wishbone_bd_ram_n20284,
         p_wishbone_bd_ram_n20285, p_wishbone_bd_ram_n20286,
         p_wishbone_bd_ram_n20287, p_wishbone_bd_ram_n20288,
         p_wishbone_bd_ram_n20289, p_wishbone_bd_ram_n20290,
         p_wishbone_bd_ram_n20291, p_wishbone_bd_ram_n20292,
         p_wishbone_bd_ram_n20293, p_wishbone_bd_ram_n20294,
         p_wishbone_bd_ram_n20295, p_wishbone_bd_ram_n20296,
         p_wishbone_bd_ram_n20297, p_wishbone_bd_ram_n20298,
         p_wishbone_bd_ram_n20299, p_wishbone_bd_ram_n20300,
         p_wishbone_bd_ram_n20301, p_wishbone_bd_ram_n20302,
         p_wishbone_bd_ram_n20303, p_wishbone_bd_ram_n20304,
         p_wishbone_bd_ram_n20305, p_wishbone_bd_ram_n20306,
         p_wishbone_bd_ram_n20307, p_wishbone_bd_ram_n20308,
         p_wishbone_bd_ram_n20309, p_wishbone_bd_ram_n20310,
         p_wishbone_bd_ram_n20311, p_wishbone_bd_ram_n20312,
         p_wishbone_bd_ram_n20313, p_wishbone_bd_ram_n20314,
         p_wishbone_bd_ram_n20315, p_wishbone_bd_ram_n20316,
         p_wishbone_bd_ram_n20317, p_wishbone_bd_ram_n20318,
         p_wishbone_bd_ram_n20319, p_wishbone_bd_ram_n20320,
         p_wishbone_bd_ram_n20321, p_wishbone_bd_ram_n20322,
         p_wishbone_bd_ram_n20323, p_wishbone_bd_ram_n20324,
         p_wishbone_bd_ram_n20325, p_wishbone_bd_ram_n20326,
         p_wishbone_bd_ram_n20327, p_wishbone_bd_ram_n20328,
         p_wishbone_bd_ram_n20329, p_wishbone_bd_ram_n20330,
         p_wishbone_bd_ram_n20331, p_wishbone_bd_ram_n20332,
         p_wishbone_bd_ram_n20333, p_wishbone_bd_ram_n20334,
         p_wishbone_bd_ram_n20335, p_wishbone_bd_ram_n20336,
         p_wishbone_bd_ram_n20337, p_wishbone_bd_ram_n20338,
         p_wishbone_bd_ram_n20339, p_wishbone_bd_ram_n20340,
         p_wishbone_bd_ram_n20341, p_wishbone_bd_ram_n20342,
         p_wishbone_bd_ram_n20343, p_wishbone_bd_ram_n20344,
         p_wishbone_bd_ram_n20345, p_wishbone_bd_ram_n20346,
         p_wishbone_bd_ram_n20347, p_wishbone_bd_ram_n20348,
         p_wishbone_bd_ram_n20349, p_wishbone_bd_ram_n20350,
         p_wishbone_bd_ram_n20351, p_wishbone_bd_ram_n20352,
         p_wishbone_bd_ram_n20353, p_wishbone_bd_ram_n20354,
         p_wishbone_bd_ram_n20355, p_wishbone_bd_ram_n20356,
         p_wishbone_bd_ram_n20357, p_wishbone_bd_ram_n20358,
         p_wishbone_bd_ram_n20359, p_wishbone_bd_ram_n20360,
         p_wishbone_bd_ram_n20361, p_wishbone_bd_ram_n20362,
         p_wishbone_bd_ram_n20363, p_wishbone_bd_ram_n20364,
         p_wishbone_bd_ram_n20365, p_wishbone_bd_ram_n20366,
         p_wishbone_bd_ram_n20367, p_wishbone_bd_ram_n20368,
         p_wishbone_bd_ram_n20369, p_wishbone_bd_ram_n20370,
         p_wishbone_bd_ram_n20371, p_wishbone_bd_ram_n20372,
         p_wishbone_bd_ram_n20373, p_wishbone_bd_ram_n20374,
         p_wishbone_bd_ram_n20375, p_wishbone_bd_ram_n20376,
         p_wishbone_bd_ram_n20377, p_wishbone_bd_ram_n20378,
         p_wishbone_bd_ram_n20379, p_wishbone_bd_ram_n20380,
         p_wishbone_bd_ram_n20381, p_wishbone_bd_ram_n20382,
         p_wishbone_bd_ram_n20383, p_wishbone_bd_ram_n20384,
         p_wishbone_bd_ram_n20385, p_wishbone_bd_ram_n20386,
         p_wishbone_bd_ram_n20387, p_wishbone_bd_ram_n20388,
         p_wishbone_bd_ram_n20389, p_wishbone_bd_ram_n20390,
         p_wishbone_bd_ram_n20391, p_wishbone_bd_ram_n20392,
         p_wishbone_bd_ram_n20393, p_wishbone_bd_ram_n20394,
         p_wishbone_bd_ram_n20395, p_wishbone_bd_ram_n20396,
         p_wishbone_bd_ram_n20397, p_wishbone_bd_ram_n20398,
         p_wishbone_bd_ram_n20399, p_wishbone_bd_ram_n20400,
         p_wishbone_bd_ram_n20401, p_wishbone_bd_ram_n20402,
         p_wishbone_bd_ram_n20403, p_wishbone_bd_ram_n20404,
         p_wishbone_bd_ram_n20405, p_wishbone_bd_ram_n20406,
         p_wishbone_bd_ram_n20407, p_wishbone_bd_ram_n20408,
         p_wishbone_bd_ram_n20409, p_wishbone_bd_ram_n20410,
         p_wishbone_bd_ram_n20411, p_wishbone_bd_ram_n20412,
         p_wishbone_bd_ram_n20413, p_wishbone_bd_ram_n20414,
         p_wishbone_bd_ram_n20415, p_wishbone_bd_ram_n20416,
         p_wishbone_bd_ram_n20417, p_wishbone_bd_ram_n20418,
         p_wishbone_bd_ram_n20419, p_wishbone_bd_ram_n20420,
         p_wishbone_bd_ram_n20421, p_wishbone_bd_ram_n20422,
         p_wishbone_bd_ram_n20423, p_wishbone_bd_ram_n20424,
         p_wishbone_bd_ram_n20425, p_wishbone_bd_ram_n20426,
         p_wishbone_bd_ram_n20427, p_wishbone_bd_ram_n20428,
         p_wishbone_bd_ram_n20429, p_wishbone_bd_ram_n20430,
         p_wishbone_bd_ram_n20431, p_wishbone_bd_ram_n20432,
         p_wishbone_bd_ram_n20433, p_wishbone_bd_ram_n20434,
         p_wishbone_bd_ram_n20435, p_wishbone_bd_ram_n20436,
         p_wishbone_bd_ram_n20437, p_wishbone_bd_ram_n20438,
         p_wishbone_bd_ram_n20439, p_wishbone_bd_ram_n20440,
         p_wishbone_bd_ram_n20441, p_wishbone_bd_ram_n20442,
         p_wishbone_bd_ram_n20443, p_wishbone_bd_ram_n20444,
         p_wishbone_bd_ram_n20445, p_wishbone_bd_ram_n20446,
         p_wishbone_bd_ram_n20447, p_wishbone_bd_ram_n20448,
         p_wishbone_bd_ram_n20449, p_wishbone_bd_ram_n20450,
         p_wishbone_bd_ram_n20451, p_wishbone_bd_ram_n20452,
         p_wishbone_bd_ram_n20453, p_wishbone_bd_ram_n20454,
         p_wishbone_bd_ram_n20455, p_wishbone_bd_ram_n20456,
         p_wishbone_bd_ram_n20457, p_wishbone_bd_ram_n20458,
         p_wishbone_bd_ram_n20459, p_wishbone_bd_ram_n20460,
         p_wishbone_bd_ram_n20461, p_wishbone_bd_ram_n20462,
         p_wishbone_bd_ram_n20463, p_wishbone_bd_ram_n20464,
         p_wishbone_bd_ram_n20465, p_wishbone_bd_ram_n20466,
         p_wishbone_bd_ram_n20467, p_wishbone_bd_ram_n20468,
         p_wishbone_bd_ram_n20469, p_wishbone_bd_ram_n20470,
         p_wishbone_bd_ram_n20471, p_wishbone_bd_ram_n20472,
         p_wishbone_bd_ram_n20473, p_wishbone_bd_ram_n20474,
         p_wishbone_bd_ram_n20475, p_wishbone_bd_ram_n20476,
         p_wishbone_bd_ram_n20477, p_wishbone_bd_ram_n20478,
         p_wishbone_bd_ram_n20479, p_wishbone_bd_ram_n20480,
         p_wishbone_bd_ram_n20481, p_wishbone_bd_ram_n20482,
         p_wishbone_bd_ram_n20483, p_wishbone_bd_ram_n20484,
         p_wishbone_bd_ram_n20485, p_wishbone_bd_ram_n20486,
         p_wishbone_bd_ram_n20487, p_wishbone_bd_ram_n20488,
         p_wishbone_bd_ram_n20489, p_wishbone_bd_ram_n20490,
         p_wishbone_bd_ram_n20491, p_wishbone_bd_ram_n20492,
         p_wishbone_bd_ram_n20493, p_wishbone_bd_ram_n20494,
         p_wishbone_bd_ram_n20495, p_wishbone_bd_ram_n20496,
         p_wishbone_bd_ram_n20497, p_wishbone_bd_ram_n20498,
         p_wishbone_bd_ram_n20499, p_wishbone_bd_ram_n20500,
         p_wishbone_bd_ram_n20501, p_wishbone_bd_ram_n20502,
         p_wishbone_bd_ram_n20503, p_wishbone_bd_ram_n20504,
         p_wishbone_bd_ram_n20505, p_wishbone_bd_ram_n20506,
         p_wishbone_bd_ram_n20507, p_wishbone_bd_ram_n20508,
         p_wishbone_bd_ram_n20509, p_wishbone_bd_ram_n20510,
         p_wishbone_bd_ram_n20511, p_wishbone_bd_ram_n20512,
         p_wishbone_bd_ram_n20513, p_wishbone_bd_ram_n20514,
         p_wishbone_bd_ram_n20515, p_wishbone_bd_ram_n20516,
         p_wishbone_bd_ram_n20517, p_wishbone_bd_ram_n20518,
         p_wishbone_bd_ram_n20519, p_wishbone_bd_ram_n20520,
         p_wishbone_bd_ram_n20521, p_wishbone_bd_ram_n20522,
         p_wishbone_bd_ram_n20523, p_wishbone_bd_ram_n20524,
         p_wishbone_bd_ram_n20525, p_wishbone_bd_ram_n20526,
         p_wishbone_bd_ram_n20527, p_wishbone_bd_ram_n20528,
         p_wishbone_bd_ram_n20529, p_wishbone_bd_ram_n20530,
         p_wishbone_bd_ram_n20531, p_wishbone_bd_ram_n20532,
         p_wishbone_bd_ram_n20533, p_wishbone_bd_ram_n20534,
         p_wishbone_bd_ram_n20535, p_wishbone_bd_ram_n20536,
         p_wishbone_bd_ram_n20537, p_wishbone_bd_ram_n20538,
         p_wishbone_bd_ram_n20539, p_wishbone_bd_ram_n20540,
         p_wishbone_bd_ram_n20541, p_wishbone_bd_ram_n20542,
         p_wishbone_bd_ram_n20543, p_wishbone_bd_ram_n20544,
         p_wishbone_bd_ram_n20545, p_wishbone_bd_ram_n20546,
         p_wishbone_bd_ram_n20547, p_wishbone_bd_ram_n20548,
         p_wishbone_bd_ram_n20549, p_wishbone_bd_ram_n20550,
         p_wishbone_bd_ram_n20551, p_wishbone_bd_ram_n20552,
         p_wishbone_bd_ram_n20553, p_wishbone_bd_ram_n20554,
         p_wishbone_bd_ram_n20555, p_wishbone_bd_ram_n20556,
         p_wishbone_bd_ram_n20557, p_wishbone_bd_ram_n20558,
         p_wishbone_bd_ram_n20559, p_wishbone_bd_ram_n20560,
         p_wishbone_bd_ram_n20561, p_wishbone_bd_ram_n20562,
         p_wishbone_bd_ram_n20563, p_wishbone_bd_ram_n20564,
         p_wishbone_bd_ram_n20565, p_wishbone_bd_ram_n20566,
         p_wishbone_bd_ram_n20567, p_wishbone_bd_ram_n20568,
         p_wishbone_bd_ram_n20569, p_wishbone_bd_ram_n20570,
         p_wishbone_bd_ram_n20571, p_wishbone_bd_ram_n20572,
         p_wishbone_bd_ram_n20573, p_wishbone_bd_ram_n20574,
         p_wishbone_bd_ram_n20575, p_wishbone_bd_ram_n20576,
         p_wishbone_bd_ram_n20577, p_wishbone_bd_ram_n20578,
         p_wishbone_bd_ram_n20579, p_wishbone_bd_ram_n20580,
         p_wishbone_bd_ram_n20581, p_wishbone_bd_ram_n20582,
         p_wishbone_bd_ram_n20583, p_wishbone_bd_ram_n20584,
         p_wishbone_bd_ram_n20585, p_wishbone_bd_ram_n20586,
         p_wishbone_bd_ram_n20587, p_wishbone_bd_ram_n20588,
         p_wishbone_bd_ram_n20589, p_wishbone_bd_ram_n20590,
         p_wishbone_bd_ram_n20591, p_wishbone_bd_ram_n20592,
         p_wishbone_bd_ram_n20593, p_wishbone_bd_ram_n20594,
         p_wishbone_bd_ram_n20595, p_wishbone_bd_ram_n20596,
         p_wishbone_bd_ram_n20597, p_wishbone_bd_ram_n20598,
         p_wishbone_bd_ram_n20599, p_wishbone_bd_ram_n20600,
         p_wishbone_bd_ram_n20601, p_wishbone_bd_ram_n20602,
         p_wishbone_bd_ram_n20603, p_wishbone_bd_ram_n20604,
         p_wishbone_bd_ram_n20605, p_wishbone_bd_ram_n20606,
         p_wishbone_bd_ram_n20607, p_wishbone_bd_ram_n20608,
         p_wishbone_bd_ram_n20609, p_wishbone_bd_ram_n20610,
         p_wishbone_bd_ram_n20611, p_wishbone_bd_ram_n20612,
         p_wishbone_bd_ram_n20613, p_wishbone_bd_ram_n20614,
         p_wishbone_bd_ram_n20615, p_wishbone_bd_ram_n20616,
         p_wishbone_bd_ram_n20617, p_wishbone_bd_ram_n20618,
         p_wishbone_bd_ram_n20619, p_wishbone_bd_ram_n20620,
         p_wishbone_bd_ram_n20621, p_wishbone_bd_ram_n20622,
         p_wishbone_bd_ram_n20623, p_wishbone_bd_ram_n20624,
         p_wishbone_bd_ram_n20625, p_wishbone_bd_ram_n20626,
         p_wishbone_bd_ram_n20627, p_wishbone_bd_ram_n20628,
         p_wishbone_bd_ram_n20629, p_wishbone_bd_ram_n20630,
         p_wishbone_bd_ram_n20631, p_wishbone_bd_ram_n20632,
         p_wishbone_bd_ram_n20633, p_wishbone_bd_ram_n20634,
         p_wishbone_bd_ram_n20635, p_wishbone_bd_ram_n20636,
         p_wishbone_bd_ram_n20637, p_wishbone_bd_ram_n20638,
         p_wishbone_bd_ram_n20639, p_wishbone_bd_ram_n20640,
         p_wishbone_bd_ram_n20641, p_wishbone_bd_ram_n20642,
         p_wishbone_bd_ram_n20643, p_wishbone_bd_ram_n20644,
         p_wishbone_bd_ram_n20645, p_wishbone_bd_ram_n20646,
         p_wishbone_bd_ram_n20647, p_wishbone_bd_ram_n20648,
         p_wishbone_bd_ram_n20649, p_wishbone_bd_ram_n20650,
         p_wishbone_bd_ram_n20651, p_wishbone_bd_ram_n20652,
         p_wishbone_bd_ram_n20653, p_wishbone_bd_ram_n20654,
         p_wishbone_bd_ram_n20655, p_wishbone_bd_ram_n20656,
         p_wishbone_bd_ram_n20657, p_wishbone_bd_ram_n20658,
         p_wishbone_bd_ram_n20659, p_wishbone_bd_ram_n20660,
         p_wishbone_bd_ram_n20661, p_wishbone_bd_ram_n20662,
         p_wishbone_bd_ram_n20663, p_wishbone_bd_ram_n20664,
         p_wishbone_bd_ram_n20665, p_wishbone_bd_ram_n20666,
         p_wishbone_bd_ram_n20667, p_wishbone_bd_ram_n20668,
         p_wishbone_bd_ram_n20669, p_wishbone_bd_ram_n20670,
         p_wishbone_bd_ram_n20671, p_wishbone_bd_ram_n20672,
         p_wishbone_bd_ram_n20673, p_wishbone_bd_ram_n20674,
         p_wishbone_bd_ram_n20675, p_wishbone_bd_ram_n20676,
         p_wishbone_bd_ram_n20677, p_wishbone_bd_ram_n20678,
         p_wishbone_bd_ram_n20679, p_wishbone_bd_ram_n20680,
         p_wishbone_bd_ram_n20681, p_wishbone_bd_ram_n20682,
         p_wishbone_bd_ram_n20683, p_wishbone_bd_ram_n20684,
         p_wishbone_bd_ram_n20685, p_wishbone_bd_ram_n20686,
         p_wishbone_bd_ram_n20687, p_wishbone_bd_ram_n20688,
         p_wishbone_bd_ram_n20689, p_wishbone_bd_ram_n20690,
         p_wishbone_bd_ram_n20691, p_wishbone_bd_ram_n20692,
         p_wishbone_bd_ram_n20693, p_wishbone_bd_ram_n20694,
         p_wishbone_bd_ram_n20695, p_wishbone_bd_ram_n20696,
         p_wishbone_bd_ram_n20697, p_wishbone_bd_ram_n20698,
         p_wishbone_bd_ram_n20699, p_wishbone_bd_ram_n20700,
         p_wishbone_bd_ram_n20701, p_wishbone_bd_ram_n20702,
         p_wishbone_bd_ram_n20703, p_wishbone_bd_ram_n20704,
         p_wishbone_bd_ram_n20705, p_wishbone_bd_ram_n20706,
         p_wishbone_bd_ram_n20707, p_wishbone_bd_ram_n20708,
         p_wishbone_bd_ram_n20709, p_wishbone_bd_ram_n20710,
         p_wishbone_bd_ram_n20711, p_wishbone_bd_ram_n20712,
         p_wishbone_bd_ram_n20713, p_wishbone_bd_ram_n20714,
         p_wishbone_bd_ram_n20715, p_wishbone_bd_ram_n20716,
         p_wishbone_bd_ram_n20717, p_wishbone_bd_ram_n20718,
         p_wishbone_bd_ram_n20719, p_wishbone_bd_ram_n20720,
         p_wishbone_bd_ram_n20721, p_wishbone_bd_ram_n20722,
         p_wishbone_bd_ram_n20723, p_wishbone_bd_ram_n20724,
         p_wishbone_bd_ram_n20725, p_wishbone_bd_ram_n20726,
         p_wishbone_bd_ram_n20727, p_wishbone_bd_ram_n20728,
         p_wishbone_bd_ram_n20729, p_wishbone_bd_ram_n20730,
         p_wishbone_bd_ram_n20731, p_wishbone_bd_ram_n20732,
         p_wishbone_bd_ram_n20733, p_wishbone_bd_ram_n20734,
         p_wishbone_bd_ram_n20735, p_wishbone_bd_ram_n20736,
         p_wishbone_bd_ram_n20737, p_wishbone_bd_ram_n20738,
         p_wishbone_bd_ram_n20739, p_wishbone_bd_ram_n20740,
         p_wishbone_bd_ram_n20741, p_wishbone_bd_ram_n20742,
         p_wishbone_bd_ram_n20743, p_wishbone_bd_ram_n20744,
         p_wishbone_bd_ram_n20745, p_wishbone_bd_ram_n20746,
         p_wishbone_bd_ram_n20747, p_wishbone_bd_ram_n20748,
         p_wishbone_bd_ram_n20749, p_wishbone_bd_ram_n20750,
         p_wishbone_bd_ram_n20751, p_wishbone_bd_ram_n20752,
         p_wishbone_bd_ram_n20753, p_wishbone_bd_ram_n20754,
         p_wishbone_bd_ram_n20755, p_wishbone_bd_ram_n20756,
         p_wishbone_bd_ram_n20757, p_wishbone_bd_ram_n20758,
         p_wishbone_bd_ram_n20759, p_wishbone_bd_ram_n20760,
         p_wishbone_bd_ram_n20761, p_wishbone_bd_ram_n20762,
         p_wishbone_bd_ram_n20763, p_wishbone_bd_ram_n20764,
         p_wishbone_bd_ram_n20765, p_wishbone_bd_ram_n20766,
         p_wishbone_bd_ram_n20767, p_wishbone_bd_ram_n20768,
         p_wishbone_bd_ram_n20769, p_wishbone_bd_ram_n20770,
         p_wishbone_bd_ram_n20771, p_wishbone_bd_ram_n20772,
         p_wishbone_bd_ram_n20773, p_wishbone_bd_ram_n20774,
         p_wishbone_bd_ram_n20775, p_wishbone_bd_ram_n20776,
         p_wishbone_bd_ram_n20777, p_wishbone_bd_ram_n20778,
         p_wishbone_bd_ram_n20779, p_wishbone_bd_ram_n20780,
         p_wishbone_bd_ram_n20781, p_wishbone_bd_ram_n20782,
         p_wishbone_bd_ram_n20783, p_wishbone_bd_ram_n20784,
         p_wishbone_bd_ram_n20785, p_wishbone_bd_ram_n20786,
         p_wishbone_bd_ram_n20787, p_wishbone_bd_ram_n20788,
         p_wishbone_bd_ram_n20789, p_wishbone_bd_ram_n20790,
         p_wishbone_bd_ram_n20791, p_wishbone_bd_ram_n20792,
         p_wishbone_bd_ram_n20793, p_wishbone_bd_ram_n20794,
         p_wishbone_bd_ram_n20795, p_wishbone_bd_ram_n20796,
         p_wishbone_bd_ram_n20797, p_wishbone_bd_ram_n20798,
         p_wishbone_bd_ram_n20799, p_wishbone_bd_ram_n20800,
         p_wishbone_bd_ram_n20801, p_wishbone_bd_ram_n20802,
         p_wishbone_bd_ram_n20803, p_wishbone_bd_ram_n20804,
         p_wishbone_bd_ram_n20805, p_wishbone_bd_ram_n20806,
         p_wishbone_bd_ram_n20807, p_wishbone_bd_ram_n20808,
         p_wishbone_bd_ram_n20809, p_wishbone_bd_ram_n20810,
         p_wishbone_bd_ram_n20811, p_wishbone_bd_ram_n20812,
         p_wishbone_bd_ram_n20813, p_wishbone_bd_ram_n20814,
         p_wishbone_bd_ram_n20815, p_wishbone_bd_ram_n20816,
         p_wishbone_bd_ram_n20817, p_wishbone_bd_ram_n20818,
         p_wishbone_bd_ram_n20819, p_wishbone_bd_ram_n20820,
         p_wishbone_bd_ram_n20821, p_wishbone_bd_ram_n20822,
         p_wishbone_bd_ram_n20823, p_wishbone_bd_ram_n20824,
         p_wishbone_bd_ram_n20825, p_wishbone_bd_ram_n20826,
         p_wishbone_bd_ram_n20827, p_wishbone_bd_ram_n20828,
         p_wishbone_bd_ram_n20829, p_wishbone_bd_ram_n20830,
         p_wishbone_bd_ram_n20831, p_wishbone_bd_ram_n20832,
         p_wishbone_bd_ram_n20833, p_wishbone_bd_ram_n20834,
         p_wishbone_bd_ram_n20835, p_wishbone_bd_ram_n20836,
         p_wishbone_bd_ram_n20837, p_wishbone_bd_ram_n20838,
         p_wishbone_bd_ram_n20839, p_wishbone_bd_ram_n20840,
         p_wishbone_bd_ram_n20841, p_wishbone_bd_ram_n20842,
         p_wishbone_bd_ram_n20843, p_wishbone_bd_ram_n20844,
         p_wishbone_bd_ram_n20845, p_wishbone_bd_ram_n20846,
         p_wishbone_bd_ram_n20847, p_wishbone_bd_ram_n20848,
         p_wishbone_bd_ram_n20849, p_wishbone_bd_ram_n20850,
         p_wishbone_bd_ram_n20851, p_wishbone_bd_ram_n20852,
         p_wishbone_bd_ram_n20853, p_wishbone_bd_ram_n20854,
         p_wishbone_bd_ram_n20855, p_wishbone_bd_ram_n20856,
         p_wishbone_bd_ram_n20857, p_wishbone_bd_ram_n20858,
         p_wishbone_bd_ram_n20859, p_wishbone_bd_ram_n20860,
         p_wishbone_bd_ram_n20861, p_wishbone_bd_ram_n20862,
         p_wishbone_bd_ram_n20863, p_wishbone_bd_ram_n20864,
         p_wishbone_bd_ram_n20865, p_wishbone_bd_ram_n20866,
         p_wishbone_bd_ram_n20867, p_wishbone_bd_ram_n20868,
         p_wishbone_bd_ram_n20869, p_wishbone_bd_ram_n20870,
         p_wishbone_bd_ram_n20871, p_wishbone_bd_ram_n20872,
         p_wishbone_bd_ram_n20873, p_wishbone_bd_ram_n20874,
         p_wishbone_bd_ram_n20875, p_wishbone_bd_ram_n20876,
         p_wishbone_bd_ram_n20877, p_wishbone_bd_ram_n20878,
         p_wishbone_bd_ram_n20879, p_wishbone_bd_ram_n20880,
         p_wishbone_bd_ram_n20881, p_wishbone_bd_ram_n20882,
         p_wishbone_bd_ram_n20883, p_wishbone_bd_ram_n20884,
         p_wishbone_bd_ram_n20885, p_wishbone_bd_ram_n20886,
         p_wishbone_bd_ram_n20887, p_wishbone_bd_ram_n20888,
         p_wishbone_bd_ram_n20889, p_wishbone_bd_ram_n20890,
         p_wishbone_bd_ram_n20891, p_wishbone_bd_ram_n20892,
         p_wishbone_bd_ram_n20893, p_wishbone_bd_ram_n20894,
         p_wishbone_bd_ram_n20895, p_wishbone_bd_ram_n20896,
         p_wishbone_bd_ram_n20897, p_wishbone_bd_ram_n20898,
         p_wishbone_bd_ram_n20899, p_wishbone_bd_ram_n20900,
         p_wishbone_bd_ram_n20901, p_wishbone_bd_ram_n20902,
         p_wishbone_bd_ram_n20903, p_wishbone_bd_ram_n20904,
         p_wishbone_bd_ram_n20905, p_wishbone_bd_ram_n20906,
         p_wishbone_bd_ram_n20907, p_wishbone_bd_ram_n20908,
         p_wishbone_bd_ram_n20909, p_wishbone_bd_ram_n20910,
         p_wishbone_bd_ram_n20911, p_wishbone_bd_ram_n20912,
         p_wishbone_bd_ram_n20913, p_wishbone_bd_ram_n20914,
         p_wishbone_bd_ram_n20915, p_wishbone_bd_ram_n20916,
         p_wishbone_bd_ram_n20917, p_wishbone_bd_ram_n20918,
         p_wishbone_bd_ram_n20919, p_wishbone_bd_ram_n20920,
         p_wishbone_bd_ram_n20921, p_wishbone_bd_ram_n20922,
         p_wishbone_bd_ram_n20923, p_wishbone_bd_ram_n20924,
         p_wishbone_bd_ram_n20925, p_wishbone_bd_ram_n20926,
         p_wishbone_bd_ram_n20927, p_wishbone_bd_ram_n20928,
         p_wishbone_bd_ram_n20929, p_wishbone_bd_ram_n20930,
         p_wishbone_bd_ram_n20931, p_wishbone_bd_ram_n20932,
         p_wishbone_bd_ram_n20933, p_wishbone_bd_ram_n20934,
         p_wishbone_bd_ram_n20935, p_wishbone_bd_ram_n20936,
         p_wishbone_bd_ram_n20937, p_wishbone_bd_ram_n20938,
         p_wishbone_bd_ram_n20939, p_wishbone_bd_ram_n20940,
         p_wishbone_bd_ram_n20941, p_wishbone_bd_ram_n20942,
         p_wishbone_bd_ram_n20943, p_wishbone_bd_ram_n20944,
         p_wishbone_bd_ram_n20945, p_wishbone_bd_ram_n20946,
         p_wishbone_bd_ram_n20947, p_wishbone_bd_ram_n20948,
         p_wishbone_bd_ram_n20949, p_wishbone_bd_ram_n20950,
         p_wishbone_bd_ram_n20951, p_wishbone_bd_ram_n20952,
         p_wishbone_bd_ram_n20953, p_wishbone_bd_ram_n20954,
         p_wishbone_bd_ram_n20955, p_wishbone_bd_ram_n20956,
         p_wishbone_bd_ram_n20957, p_wishbone_bd_ram_n20958,
         p_wishbone_bd_ram_n20959, p_wishbone_bd_ram_n20960,
         p_wishbone_bd_ram_n20961, p_wishbone_bd_ram_n20962,
         p_wishbone_bd_ram_n20963, p_wishbone_bd_ram_n20964,
         p_wishbone_bd_ram_n20965, p_wishbone_bd_ram_n20966,
         p_wishbone_bd_ram_n20967, p_wishbone_bd_ram_n20968,
         p_wishbone_bd_ram_n20969, p_wishbone_bd_ram_n20970,
         p_wishbone_bd_ram_n20971, p_wishbone_bd_ram_n20972,
         p_wishbone_bd_ram_n20973, p_wishbone_bd_ram_n20974,
         p_wishbone_bd_ram_n20975, p_wishbone_bd_ram_n20976,
         p_wishbone_bd_ram_n20977, p_wishbone_bd_ram_n20978,
         p_wishbone_bd_ram_n20979, p_wishbone_bd_ram_n20980,
         p_wishbone_bd_ram_n20981, p_wishbone_bd_ram_n20982,
         p_wishbone_bd_ram_n20983, p_wishbone_bd_ram_n20984,
         p_wishbone_bd_ram_n20985, p_wishbone_bd_ram_n20986,
         p_wishbone_bd_ram_n20987, p_wishbone_bd_ram_n20988,
         p_wishbone_bd_ram_n20989, p_wishbone_bd_ram_n20990,
         p_wishbone_bd_ram_n20991, p_wishbone_bd_ram_n20992,
         p_wishbone_bd_ram_n20993, p_wishbone_bd_ram_n20994,
         p_wishbone_bd_ram_n20995, p_wishbone_bd_ram_n20996,
         p_wishbone_bd_ram_n20997, p_wishbone_bd_ram_n20998,
         p_wishbone_bd_ram_n20999, p_wishbone_bd_ram_n21000,
         p_wishbone_bd_ram_n21001, p_wishbone_bd_ram_n21002,
         p_wishbone_bd_ram_n21003, p_wishbone_bd_ram_n21004,
         p_wishbone_bd_ram_n21005, p_wishbone_bd_ram_n21006,
         p_wishbone_bd_ram_n21007, p_wishbone_bd_ram_n21008,
         p_wishbone_bd_ram_n21009, p_wishbone_bd_ram_n21010,
         p_wishbone_bd_ram_n21011, p_wishbone_bd_ram_n21012,
         p_wishbone_bd_ram_n21013, p_wishbone_bd_ram_n21014,
         p_wishbone_bd_ram_n21015, p_wishbone_bd_ram_n21016,
         p_wishbone_bd_ram_n21017, p_wishbone_bd_ram_n21018,
         p_wishbone_bd_ram_n21019, p_wishbone_bd_ram_n21020,
         p_wishbone_bd_ram_n21021, p_wishbone_bd_ram_n21022,
         p_wishbone_bd_ram_n21023, p_wishbone_bd_ram_n21024,
         p_wishbone_bd_ram_n21025, p_wishbone_bd_ram_n21026,
         p_wishbone_bd_ram_n21027, p_wishbone_bd_ram_n21028,
         p_wishbone_bd_ram_n21029, p_wishbone_bd_ram_n21030,
         p_wishbone_bd_ram_n21031, p_wishbone_bd_ram_n21032,
         p_wishbone_bd_ram_n21033, p_wishbone_bd_ram_n21034,
         p_wishbone_bd_ram_n21035, p_wishbone_bd_ram_n21036,
         p_wishbone_bd_ram_n21037, p_wishbone_bd_ram_n21038,
         p_wishbone_bd_ram_n21039, p_wishbone_bd_ram_n21040,
         p_wishbone_bd_ram_n21041, p_wishbone_bd_ram_n21042,
         p_wishbone_bd_ram_n21043, p_wishbone_bd_ram_n21044,
         p_wishbone_bd_ram_n21045, p_wishbone_bd_ram_n21046,
         p_wishbone_bd_ram_n21047, p_wishbone_bd_ram_n21048,
         p_wishbone_bd_ram_n21049, p_wishbone_bd_ram_n21050,
         p_wishbone_bd_ram_n21051, p_wishbone_bd_ram_n21052,
         p_wishbone_bd_ram_n21053, p_wishbone_bd_ram_n21054,
         p_wishbone_bd_ram_n21055, p_wishbone_bd_ram_n21056,
         p_wishbone_bd_ram_n21057, p_wishbone_bd_ram_n21058,
         p_wishbone_bd_ram_n21059, p_wishbone_bd_ram_n21060,
         p_wishbone_bd_ram_n21061, p_wishbone_bd_ram_n21062,
         p_wishbone_bd_ram_n21063, p_wishbone_bd_ram_n21064,
         p_wishbone_bd_ram_n21065, p_wishbone_bd_ram_n21066,
         p_wishbone_bd_ram_n21067, p_wishbone_bd_ram_n21068,
         p_wishbone_bd_ram_n21069, p_wishbone_bd_ram_n21070,
         p_wishbone_bd_ram_n21071, p_wishbone_bd_ram_n21072,
         p_wishbone_bd_ram_n21073, p_wishbone_bd_ram_n21074,
         p_wishbone_bd_ram_n21075, p_wishbone_bd_ram_n21076,
         p_wishbone_bd_ram_n21077, p_wishbone_bd_ram_n21078,
         p_wishbone_bd_ram_n21079, p_wishbone_bd_ram_n21080,
         p_wishbone_bd_ram_n21081, p_wishbone_bd_ram_n21082,
         p_wishbone_bd_ram_n21083, p_wishbone_bd_ram_n21084,
         p_wishbone_bd_ram_n21085, p_wishbone_bd_ram_n21086,
         p_wishbone_bd_ram_n21087, p_wishbone_bd_ram_n21088,
         p_wishbone_bd_ram_n21089, p_wishbone_bd_ram_n21090,
         p_wishbone_bd_ram_n21091, p_wishbone_bd_ram_n21092,
         p_wishbone_bd_ram_n21093, p_wishbone_bd_ram_n21094,
         p_wishbone_bd_ram_n21095, p_wishbone_bd_ram_n21096,
         p_wishbone_bd_ram_n21097, p_wishbone_bd_ram_n21098,
         p_wishbone_bd_ram_n21099, p_wishbone_bd_ram_n21100,
         p_wishbone_bd_ram_n21101, p_wishbone_bd_ram_n21102,
         p_wishbone_bd_ram_n21103, p_wishbone_bd_ram_n21104,
         p_wishbone_bd_ram_n21105, p_wishbone_bd_ram_n21106,
         p_wishbone_bd_ram_n21107, p_wishbone_bd_ram_n21108,
         p_wishbone_bd_ram_n21109, p_wishbone_bd_ram_n21110,
         p_wishbone_bd_ram_n21111, p_wishbone_bd_ram_n21112,
         p_wishbone_bd_ram_n21113, p_wishbone_bd_ram_n21114,
         p_wishbone_bd_ram_n21115, p_wishbone_bd_ram_n21116,
         p_wishbone_bd_ram_n21117, p_wishbone_bd_ram_n21118,
         p_wishbone_bd_ram_n21119, p_wishbone_bd_ram_n21120,
         p_wishbone_bd_ram_n21121, p_wishbone_bd_ram_n21122,
         p_wishbone_bd_ram_n21123, p_wishbone_bd_ram_n21124,
         p_wishbone_bd_ram_n21125, p_wishbone_bd_ram_n21126,
         p_wishbone_bd_ram_n21127, p_wishbone_bd_ram_n21128,
         p_wishbone_bd_ram_n21129, p_wishbone_bd_ram_n21130,
         p_wishbone_bd_ram_n21131, p_wishbone_bd_ram_n21132,
         p_wishbone_bd_ram_n21133, p_wishbone_bd_ram_n21134,
         p_wishbone_bd_ram_n21135, p_wishbone_bd_ram_n21136,
         p_wishbone_bd_ram_n21137, p_wishbone_bd_ram_n21138,
         p_wishbone_bd_ram_n21139, p_wishbone_bd_ram_n21140,
         p_wishbone_bd_ram_n21141, p_wishbone_bd_ram_n21142,
         p_wishbone_bd_ram_n21143, p_wishbone_bd_ram_n21144,
         p_wishbone_bd_ram_n21145, p_wishbone_bd_ram_n21146,
         p_wishbone_bd_ram_n21147, p_wishbone_bd_ram_n21148,
         p_wishbone_bd_ram_n21149, p_wishbone_bd_ram_n21150,
         p_wishbone_bd_ram_n21151, p_wishbone_bd_ram_n21152,
         p_wishbone_bd_ram_n21153, p_wishbone_bd_ram_n21154,
         p_wishbone_bd_ram_n21155, p_wishbone_bd_ram_n21156,
         p_wishbone_bd_ram_n21157, p_wishbone_bd_ram_n21158,
         p_wishbone_bd_ram_n21159, p_wishbone_bd_ram_n21160,
         p_wishbone_bd_ram_n21161, p_wishbone_bd_ram_n21162,
         p_wishbone_bd_ram_n21163, p_wishbone_bd_ram_n21164,
         p_wishbone_bd_ram_n21165, p_wishbone_bd_ram_n21166,
         p_wishbone_bd_ram_n21167, p_wishbone_bd_ram_n21168,
         p_wishbone_bd_ram_n21169, p_wishbone_bd_ram_n21170,
         p_wishbone_bd_ram_n21171, p_wishbone_bd_ram_n21172,
         p_wishbone_bd_ram_n21173, p_wishbone_bd_ram_n21174,
         p_wishbone_bd_ram_n21175, p_wishbone_bd_ram_n21176,
         p_wishbone_bd_ram_n21177, p_wishbone_bd_ram_n21178,
         p_wishbone_bd_ram_n21179, p_wishbone_bd_ram_n21180,
         p_wishbone_bd_ram_n21181, p_wishbone_bd_ram_n21182,
         p_wishbone_bd_ram_n21183, p_wishbone_bd_ram_n21184,
         p_wishbone_bd_ram_n21185, p_wishbone_bd_ram_n21186,
         p_wishbone_bd_ram_n21187, p_wishbone_bd_ram_n21188,
         p_wishbone_bd_ram_n21189, p_wishbone_bd_ram_n21190,
         p_wishbone_bd_ram_n21191, p_wishbone_bd_ram_n21192,
         p_wishbone_bd_ram_n21193, p_wishbone_bd_ram_n21194,
         p_wishbone_bd_ram_n21195, p_wishbone_bd_ram_n21196,
         p_wishbone_bd_ram_n21197, p_wishbone_bd_ram_n21198,
         p_wishbone_bd_ram_n21199, p_wishbone_bd_ram_n21200,
         p_wishbone_bd_ram_n21201, p_wishbone_bd_ram_n21202,
         p_wishbone_bd_ram_n21203, p_wishbone_bd_ram_n21204,
         p_wishbone_bd_ram_n21205, p_wishbone_bd_ram_n21206,
         p_wishbone_bd_ram_n21207, p_wishbone_bd_ram_n21208,
         p_wishbone_bd_ram_n21209, p_wishbone_bd_ram_n21210,
         p_wishbone_bd_ram_n21211, p_wishbone_bd_ram_n21212,
         p_wishbone_bd_ram_n21213, p_wishbone_bd_ram_n21214,
         p_wishbone_bd_ram_n21215, p_wishbone_bd_ram_n21216,
         p_wishbone_bd_ram_n21217, p_wishbone_bd_ram_n21218,
         p_wishbone_bd_ram_n21219, p_wishbone_bd_ram_n21220,
         p_wishbone_bd_ram_n21221, p_wishbone_bd_ram_n21222,
         p_wishbone_bd_ram_n21223, p_wishbone_bd_ram_n21224,
         p_wishbone_bd_ram_n21225, p_wishbone_bd_ram_n21226,
         p_wishbone_bd_ram_n21227, p_wishbone_bd_ram_n21228,
         p_wishbone_bd_ram_n21229, p_wishbone_bd_ram_n21230,
         p_wishbone_bd_ram_n21231, p_wishbone_bd_ram_n21232,
         p_wishbone_bd_ram_n21233, p_wishbone_bd_ram_n21234,
         p_wishbone_bd_ram_n21235, p_wishbone_bd_ram_n21236,
         p_wishbone_bd_ram_n21237, p_wishbone_bd_ram_n21238,
         p_wishbone_bd_ram_n21239, p_wishbone_bd_ram_n21240,
         p_wishbone_bd_ram_n21241, p_wishbone_bd_ram_n21242,
         p_wishbone_bd_ram_n21243, p_wishbone_bd_ram_n21244,
         p_wishbone_bd_ram_n21245, p_wishbone_bd_ram_n21246,
         p_wishbone_bd_ram_n21247, p_wishbone_bd_ram_n21248,
         p_wishbone_bd_ram_n21249, p_wishbone_bd_ram_n21250,
         p_wishbone_bd_ram_n21251, p_wishbone_bd_ram_n21252,
         p_wishbone_bd_ram_n21253, p_wishbone_bd_ram_n21254,
         p_wishbone_bd_ram_n21255, p_wishbone_bd_ram_n21256,
         p_wishbone_bd_ram_n21257, p_wishbone_bd_ram_n21258,
         p_wishbone_bd_ram_n21259, p_wishbone_bd_ram_n21260,
         p_wishbone_bd_ram_n21261, p_wishbone_bd_ram_n21262,
         p_wishbone_bd_ram_n21263, p_wishbone_bd_ram_n21264,
         p_wishbone_bd_ram_n21265, p_wishbone_bd_ram_n21266,
         p_wishbone_bd_ram_n21267, p_wishbone_bd_ram_n21268,
         p_wishbone_bd_ram_n21269, p_wishbone_bd_ram_n21270,
         p_wishbone_bd_ram_n21271, p_wishbone_bd_ram_n21272,
         p_wishbone_bd_ram_n21273, p_wishbone_bd_ram_n21274,
         p_wishbone_bd_ram_n21275, p_wishbone_bd_ram_n21276,
         p_wishbone_bd_ram_n21277, p_wishbone_bd_ram_n21278,
         p_wishbone_bd_ram_n21279, p_wishbone_bd_ram_n21280,
         p_wishbone_bd_ram_n21281, p_wishbone_bd_ram_n21282,
         p_wishbone_bd_ram_n21283, p_wishbone_bd_ram_n21284,
         p_wishbone_bd_ram_n21285, p_wishbone_bd_ram_n21286,
         p_wishbone_bd_ram_n21287, p_wishbone_bd_ram_n21288,
         p_wishbone_bd_ram_n21289, p_wishbone_bd_ram_n21290,
         p_wishbone_bd_ram_n21291, p_wishbone_bd_ram_n21292,
         p_wishbone_bd_ram_n21293, p_wishbone_bd_ram_n21294,
         p_wishbone_bd_ram_n21295, p_wishbone_bd_ram_n21296,
         p_wishbone_bd_ram_n21297, p_wishbone_bd_ram_n21298,
         p_wishbone_bd_ram_n21299, p_wishbone_bd_ram_n21300,
         p_wishbone_bd_ram_n21301, p_wishbone_bd_ram_n21302,
         p_wishbone_bd_ram_n21303, p_wishbone_bd_ram_n21304,
         p_wishbone_bd_ram_n21305, p_wishbone_bd_ram_n21306,
         p_wishbone_bd_ram_n21307, p_wishbone_bd_ram_n21308,
         p_wishbone_bd_ram_n21309, p_wishbone_bd_ram_n21310,
         p_wishbone_bd_ram_n21311, p_wishbone_bd_ram_n21312,
         p_wishbone_bd_ram_n21313, p_wishbone_bd_ram_n21314,
         p_wishbone_bd_ram_n21315, p_wishbone_bd_ram_n21316,
         p_wishbone_bd_ram_n21317, p_wishbone_bd_ram_n21318,
         p_wishbone_bd_ram_n21319, p_wishbone_bd_ram_n21320,
         p_wishbone_bd_ram_n21321, p_wishbone_bd_ram_n21322,
         p_wishbone_bd_ram_n21323, p_wishbone_bd_ram_n21324,
         p_wishbone_bd_ram_n21325, p_wishbone_bd_ram_n21326,
         p_wishbone_bd_ram_n21327, p_wishbone_bd_ram_n21328,
         p_wishbone_bd_ram_n21329, p_wishbone_bd_ram_n21330,
         p_wishbone_bd_ram_n21331, p_wishbone_bd_ram_n21332,
         p_wishbone_bd_ram_n21333, p_wishbone_bd_ram_n21334,
         p_wishbone_bd_ram_n21335, p_wishbone_bd_ram_n21336,
         p_wishbone_bd_ram_n21337, p_wishbone_bd_ram_n21338,
         p_wishbone_bd_ram_n21339, p_wishbone_bd_ram_n21340,
         p_wishbone_bd_ram_n21341, p_wishbone_bd_ram_n21342,
         p_wishbone_bd_ram_n21343, p_wishbone_bd_ram_n21344,
         p_wishbone_bd_ram_n21345, p_wishbone_bd_ram_n21346,
         p_wishbone_bd_ram_n21347, p_wishbone_bd_ram_n21348,
         p_wishbone_bd_ram_n21349, p_wishbone_bd_ram_n21350,
         p_wishbone_bd_ram_n21351, p_wishbone_bd_ram_n21352,
         p_wishbone_bd_ram_n21353, p_wishbone_bd_ram_n21354,
         p_wishbone_bd_ram_n21355, p_wishbone_bd_ram_n21356,
         p_wishbone_bd_ram_n21357, p_wishbone_bd_ram_n21358,
         p_wishbone_bd_ram_n21359, p_wishbone_bd_ram_n21360,
         p_wishbone_bd_ram_n21361, p_wishbone_bd_ram_n21362,
         p_wishbone_bd_ram_n21363, p_wishbone_bd_ram_n21364,
         p_wishbone_bd_ram_n21365, p_wishbone_bd_ram_n21366,
         p_wishbone_bd_ram_n21367, p_wishbone_bd_ram_n21368,
         p_wishbone_bd_ram_n21369, p_wishbone_bd_ram_n21370,
         p_wishbone_bd_ram_n21371, p_wishbone_bd_ram_n21372,
         p_wishbone_bd_ram_n21373, p_wishbone_bd_ram_n21374,
         p_wishbone_bd_ram_n21375, p_wishbone_bd_ram_n21376,
         p_wishbone_bd_ram_n21377, p_wishbone_bd_ram_n21378,
         p_wishbone_bd_ram_n21379, p_wishbone_bd_ram_n21380,
         p_wishbone_bd_ram_n21381, p_wishbone_bd_ram_n21382,
         p_wishbone_bd_ram_n21383, p_wishbone_bd_ram_n21384,
         p_wishbone_bd_ram_n21385, p_wishbone_bd_ram_n21386,
         p_wishbone_bd_ram_n21387, p_wishbone_bd_ram_n21388,
         p_wishbone_bd_ram_n21389, p_wishbone_bd_ram_n21390,
         p_wishbone_bd_ram_n21391, p_wishbone_bd_ram_n21392,
         p_wishbone_bd_ram_n21393, p_wishbone_bd_ram_n21394,
         p_wishbone_bd_ram_n21395, p_wishbone_bd_ram_n21396,
         p_wishbone_bd_ram_n21397, p_wishbone_bd_ram_n21398,
         p_wishbone_bd_ram_n21399, p_wishbone_bd_ram_n21400,
         p_wishbone_bd_ram_n21401, p_wishbone_bd_ram_n21402,
         p_wishbone_bd_ram_n21403, p_wishbone_bd_ram_n21404,
         p_wishbone_bd_ram_n21405, p_wishbone_bd_ram_n21406,
         p_wishbone_bd_ram_n21407, p_wishbone_bd_ram_n21408,
         p_wishbone_bd_ram_n21409, p_wishbone_bd_ram_n21410,
         p_wishbone_bd_ram_n21411, p_wishbone_bd_ram_n21412,
         p_wishbone_bd_ram_n21413, p_wishbone_bd_ram_n21414,
         p_wishbone_bd_ram_n21415, p_wishbone_bd_ram_n21416,
         p_wishbone_bd_ram_n21417, p_wishbone_bd_ram_n21418,
         p_wishbone_bd_ram_n21419, p_wishbone_bd_ram_n21420,
         p_wishbone_bd_ram_n21421, p_wishbone_bd_ram_n21422,
         p_wishbone_bd_ram_n21423, p_wishbone_bd_ram_n21424,
         p_wishbone_bd_ram_n21425, p_wishbone_bd_ram_n21426,
         p_wishbone_bd_ram_n21427, p_wishbone_bd_ram_n21428,
         p_wishbone_bd_ram_n21429, p_wishbone_bd_ram_n21430,
         p_wishbone_bd_ram_n21431, p_wishbone_bd_ram_n21432,
         p_wishbone_bd_ram_n21433, p_wishbone_bd_ram_n21434,
         p_wishbone_bd_ram_n21435, p_wishbone_bd_ram_n21436,
         p_wishbone_bd_ram_n21437, p_wishbone_bd_ram_n21438,
         p_wishbone_bd_ram_n21439, p_wishbone_bd_ram_n21440,
         p_wishbone_bd_ram_n21441, p_wishbone_bd_ram_n21442,
         p_wishbone_bd_ram_n21443, p_wishbone_bd_ram_n21444,
         p_wishbone_bd_ram_n21445, p_wishbone_bd_ram_n21446,
         p_wishbone_bd_ram_n21447, p_wishbone_bd_ram_n21448,
         p_wishbone_bd_ram_n21449, p_wishbone_bd_ram_n21450,
         p_wishbone_bd_ram_n21451, p_wishbone_bd_ram_n21452,
         p_wishbone_bd_ram_n21453, p_wishbone_bd_ram_n21454,
         p_wishbone_bd_ram_n21455, p_wishbone_bd_ram_n21456,
         p_wishbone_bd_ram_n21457, p_wishbone_bd_ram_n21458,
         p_wishbone_bd_ram_n21459, p_wishbone_bd_ram_n21460,
         p_wishbone_bd_ram_n21461, p_wishbone_bd_ram_n21462,
         p_wishbone_bd_ram_n21463, p_wishbone_bd_ram_n21464,
         p_wishbone_bd_ram_n21465, p_wishbone_bd_ram_n21466,
         p_wishbone_bd_ram_n21467, p_wishbone_bd_ram_n21468,
         p_wishbone_bd_ram_n21469, p_wishbone_bd_ram_n21470,
         p_wishbone_bd_ram_n21471, p_wishbone_bd_ram_n21472,
         p_wishbone_bd_ram_n21473, p_wishbone_bd_ram_n21474,
         p_wishbone_bd_ram_n21475, p_wishbone_bd_ram_n21476,
         p_wishbone_bd_ram_n21477, p_wishbone_bd_ram_n21478,
         p_wishbone_bd_ram_n21479, p_wishbone_bd_ram_n21480,
         p_wishbone_bd_ram_n21481, p_wishbone_bd_ram_n21482,
         p_wishbone_bd_ram_n21483, p_wishbone_bd_ram_n21484,
         p_wishbone_bd_ram_n21485, p_wishbone_bd_ram_n21486,
         p_wishbone_bd_ram_n21487, p_wishbone_bd_ram_n21488,
         p_wishbone_bd_ram_n21489, p_wishbone_bd_ram_n21490,
         p_wishbone_bd_ram_n21491, p_wishbone_bd_ram_n21492,
         p_wishbone_bd_ram_n21493, p_wishbone_bd_ram_n21494,
         p_wishbone_bd_ram_n21495, p_wishbone_bd_ram_n21496,
         p_wishbone_bd_ram_n21497, p_wishbone_bd_ram_n21498,
         p_wishbone_bd_ram_n21499, p_wishbone_bd_ram_n21500,
         p_wishbone_bd_ram_n21501, p_wishbone_bd_ram_n21502,
         p_wishbone_bd_ram_n21503, p_wishbone_bd_ram_n21504,
         p_wishbone_bd_ram_n21505, p_wishbone_bd_ram_n21506,
         p_wishbone_bd_ram_n21507, p_wishbone_bd_ram_n21508,
         p_wishbone_bd_ram_n21509, p_wishbone_bd_ram_n21510,
         p_wishbone_bd_ram_n21511, p_wishbone_bd_ram_n21512,
         p_wishbone_bd_ram_n21513, p_wishbone_bd_ram_n21514,
         p_wishbone_bd_ram_n21515, p_wishbone_bd_ram_n21516,
         p_wishbone_bd_ram_n21517, p_wishbone_bd_ram_n21518,
         p_wishbone_bd_ram_n21519, p_wishbone_bd_ram_n21520,
         p_wishbone_bd_ram_n21521, p_wishbone_bd_ram_n21522,
         p_wishbone_bd_ram_n21523, p_wishbone_bd_ram_n21524,
         p_wishbone_bd_ram_n21525, p_wishbone_bd_ram_n21526,
         p_wishbone_bd_ram_n21527, p_wishbone_bd_ram_n21528,
         p_wishbone_bd_ram_n21529, p_wishbone_bd_ram_n21530,
         p_wishbone_bd_ram_n21531, p_wishbone_bd_ram_n21532,
         p_wishbone_bd_ram_n21533, p_wishbone_bd_ram_n21534,
         p_wishbone_bd_ram_n21535, p_wishbone_bd_ram_n21536,
         p_wishbone_bd_ram_n21537, p_wishbone_bd_ram_n21538,
         p_wishbone_bd_ram_n21539, p_wishbone_bd_ram_n21540,
         p_wishbone_bd_ram_n21541, p_wishbone_bd_ram_n21542,
         p_wishbone_bd_ram_n21543, p_wishbone_bd_ram_n21544,
         p_wishbone_bd_ram_n21545, p_wishbone_bd_ram_n21546,
         p_wishbone_bd_ram_n21547, p_wishbone_bd_ram_n21548,
         p_wishbone_bd_ram_n21549, p_wishbone_bd_ram_n21550,
         p_wishbone_bd_ram_n21551, p_wishbone_bd_ram_n21552,
         p_wishbone_bd_ram_n21553, p_wishbone_bd_ram_n21554,
         p_wishbone_bd_ram_n21555, p_wishbone_bd_ram_n21556,
         p_wishbone_bd_ram_n21557, p_wishbone_bd_ram_n21558,
         p_wishbone_bd_ram_n21559, p_wishbone_bd_ram_n21560,
         p_wishbone_bd_ram_n21561, p_wishbone_bd_ram_n21562,
         p_wishbone_bd_ram_n21563, p_wishbone_bd_ram_n21564,
         p_wishbone_bd_ram_n21565, p_wishbone_bd_ram_n21566,
         p_wishbone_bd_ram_n21567, p_wishbone_bd_ram_n21568,
         p_wishbone_bd_ram_n21569, p_wishbone_bd_ram_n21570,
         p_wishbone_bd_ram_n21571, p_wishbone_bd_ram_n21572,
         p_wishbone_bd_ram_n21573, p_wishbone_bd_ram_n21574,
         p_wishbone_bd_ram_n21575, p_wishbone_bd_ram_n21576,
         p_wishbone_bd_ram_n21577, p_wishbone_bd_ram_n21578,
         p_wishbone_bd_ram_n21579, p_wishbone_bd_ram_n21580,
         p_wishbone_bd_ram_n21581, p_wishbone_bd_ram_n21582,
         p_wishbone_bd_ram_n21583, p_wishbone_bd_ram_n21584,
         p_wishbone_bd_ram_n21585, p_wishbone_bd_ram_n21586,
         p_wishbone_bd_ram_n21587, p_wishbone_bd_ram_n21588,
         p_wishbone_bd_ram_n21589, p_wishbone_bd_ram_n21590,
         p_wishbone_bd_ram_n21591, p_wishbone_bd_ram_n21592,
         p_wishbone_bd_ram_n21593, p_wishbone_bd_ram_n21594,
         p_wishbone_bd_ram_n21595, p_wishbone_bd_ram_n21596,
         p_wishbone_bd_ram_n21597, p_wishbone_bd_ram_n21598,
         p_wishbone_bd_ram_n21599, p_wishbone_bd_ram_n21600,
         p_wishbone_bd_ram_n21601, p_wishbone_bd_ram_n21602,
         p_wishbone_bd_ram_n21603, p_wishbone_bd_ram_n21604,
         p_wishbone_bd_ram_n21605, p_wishbone_bd_ram_n21606,
         p_wishbone_bd_ram_n21607, p_wishbone_bd_ram_n21608,
         p_wishbone_bd_ram_n21609, p_wishbone_bd_ram_n21610,
         p_wishbone_bd_ram_n21611, p_wishbone_bd_ram_n21612,
         p_wishbone_bd_ram_n21613, p_wishbone_bd_ram_n21614,
         p_wishbone_bd_ram_n21615, p_wishbone_bd_ram_n21616,
         p_wishbone_bd_ram_n21617, p_wishbone_bd_ram_n21618,
         p_wishbone_bd_ram_n21619, p_wishbone_bd_ram_n21620,
         p_wishbone_bd_ram_n21621, p_wishbone_bd_ram_n21622,
         p_wishbone_bd_ram_n21623, p_wishbone_bd_ram_n21624,
         p_wishbone_bd_ram_n21625, p_wishbone_bd_ram_n21626,
         p_wishbone_bd_ram_n21627, p_wishbone_bd_ram_n21628,
         p_wishbone_bd_ram_n21629, p_wishbone_bd_ram_n21630,
         p_wishbone_bd_ram_n21631, p_wishbone_bd_ram_n21632,
         p_wishbone_bd_ram_n21633, p_wishbone_bd_ram_n21634,
         p_wishbone_bd_ram_n21635, p_wishbone_bd_ram_n21636,
         p_wishbone_bd_ram_n21637, p_wishbone_bd_ram_n21638,
         p_wishbone_bd_ram_n21639, p_wishbone_bd_ram_n21640,
         p_wishbone_bd_ram_n21641, p_wishbone_bd_ram_n21642,
         p_wishbone_bd_ram_n21643, p_wishbone_bd_ram_n21644,
         p_wishbone_bd_ram_n21645, p_wishbone_bd_ram_n21646,
         p_wishbone_bd_ram_n21647, p_wishbone_bd_ram_n21648,
         p_wishbone_bd_ram_n21649, p_wishbone_bd_ram_n21650,
         p_wishbone_bd_ram_n21651, p_wishbone_bd_ram_n21652,
         p_wishbone_bd_ram_n21653, p_wishbone_bd_ram_n21654,
         p_wishbone_bd_ram_n21655, p_wishbone_bd_ram_n21656,
         p_wishbone_bd_ram_n21657, p_wishbone_bd_ram_n21658,
         p_wishbone_bd_ram_n21659, p_wishbone_bd_ram_n21660,
         p_wishbone_bd_ram_n21661, p_wishbone_bd_ram_n21662,
         p_wishbone_bd_ram_n21663, p_wishbone_bd_ram_n21664,
         p_wishbone_bd_ram_n21665, p_wishbone_bd_ram_n21666,
         p_wishbone_bd_ram_n21667, p_wishbone_bd_ram_n21668,
         p_wishbone_bd_ram_n21669, p_wishbone_bd_ram_n21670,
         p_wishbone_bd_ram_n21671, p_wishbone_bd_ram_n21672,
         p_wishbone_bd_ram_n21673, p_wishbone_bd_ram_n21674,
         p_wishbone_bd_ram_n21675, p_wishbone_bd_ram_n21676,
         p_wishbone_bd_ram_n21677, p_wishbone_bd_ram_n21678,
         p_wishbone_bd_ram_n21679, p_wishbone_bd_ram_n21680,
         p_wishbone_bd_ram_n21681, p_wishbone_bd_ram_n21682,
         p_wishbone_bd_ram_n21683, p_wishbone_bd_ram_n21684,
         p_wishbone_bd_ram_n21685, p_wishbone_bd_ram_n21686,
         p_wishbone_bd_ram_n21687, p_wishbone_bd_ram_n21688,
         p_wishbone_bd_ram_n21689, p_wishbone_bd_ram_n21690,
         p_wishbone_bd_ram_n21691, p_wishbone_bd_ram_n21692,
         p_wishbone_bd_ram_n21693, p_wishbone_bd_ram_n21694,
         p_wishbone_bd_ram_n21695, p_wishbone_bd_ram_n21696,
         p_wishbone_bd_ram_n21697, p_wishbone_bd_ram_n21698,
         p_wishbone_bd_ram_n21699, p_wishbone_bd_ram_n21700,
         p_wishbone_bd_ram_n21701, p_wishbone_bd_ram_n21702,
         p_wishbone_bd_ram_n21703, p_wishbone_bd_ram_n21704,
         p_wishbone_bd_ram_n21705, p_wishbone_bd_ram_n21706,
         p_wishbone_bd_ram_n21707, p_wishbone_bd_ram_n21708,
         p_wishbone_bd_ram_n21709, p_wishbone_bd_ram_n21710,
         p_wishbone_bd_ram_n21711, p_wishbone_bd_ram_n21712,
         p_wishbone_bd_ram_n21713, p_wishbone_bd_ram_n21714,
         p_wishbone_bd_ram_n21715, p_wishbone_bd_ram_n21716,
         p_wishbone_bd_ram_n21717, p_wishbone_bd_ram_n21718,
         p_wishbone_bd_ram_n21719, p_wishbone_bd_ram_n21720,
         p_wishbone_bd_ram_n21721, p_wishbone_bd_ram_n21722,
         p_wishbone_bd_ram_n21723, p_wishbone_bd_ram_n21724,
         p_wishbone_bd_ram_n21725, p_wishbone_bd_ram_n21726,
         p_wishbone_bd_ram_n21727, p_wishbone_bd_ram_n21728,
         p_wishbone_bd_ram_n21729, p_wishbone_bd_ram_n21730,
         p_wishbone_bd_ram_n21731, p_wishbone_bd_ram_n21732,
         p_wishbone_bd_ram_n21733, p_wishbone_bd_ram_n21734,
         p_wishbone_bd_ram_n21735, p_wishbone_bd_ram_n21736,
         p_wishbone_bd_ram_n21737, p_wishbone_bd_ram_n21738,
         p_wishbone_bd_ram_n21739, p_wishbone_bd_ram_n21740,
         p_wishbone_bd_ram_n21741, p_wishbone_bd_ram_n21742,
         p_wishbone_bd_ram_n21743, p_wishbone_bd_ram_n21744,
         p_wishbone_bd_ram_n21745, p_wishbone_bd_ram_n21746,
         p_wishbone_bd_ram_n21747, p_wishbone_bd_ram_n21748,
         p_wishbone_bd_ram_n21749, p_wishbone_bd_ram_n21750,
         p_wishbone_bd_ram_n21751, p_wishbone_bd_ram_n21752,
         p_wishbone_bd_ram_n21753, p_wishbone_bd_ram_n21754,
         p_wishbone_bd_ram_n21755, p_wishbone_bd_ram_n21756,
         p_wishbone_bd_ram_n21757, p_wishbone_bd_ram_n21758,
         p_wishbone_bd_ram_n21759, p_wishbone_bd_ram_n21760,
         p_wishbone_bd_ram_n21761, p_wishbone_bd_ram_n21762,
         p_wishbone_bd_ram_n21763, p_wishbone_bd_ram_n21764,
         p_wishbone_bd_ram_n21765, p_wishbone_bd_ram_n21766,
         p_wishbone_bd_ram_n21767, p_wishbone_bd_ram_n21768,
         p_wishbone_bd_ram_n21769, p_wishbone_bd_ram_n21770,
         p_wishbone_bd_ram_n21771, p_wishbone_bd_ram_n21772,
         p_wishbone_bd_ram_n21773, p_wishbone_bd_ram_n21774,
         p_wishbone_bd_ram_n21775, p_wishbone_bd_ram_n21776,
         p_wishbone_bd_ram_n21777, p_wishbone_bd_ram_n21778,
         p_wishbone_bd_ram_n21779, p_wishbone_bd_ram_n21780,
         p_wishbone_bd_ram_n21781, p_wishbone_bd_ram_n21782,
         p_wishbone_bd_ram_n21783, p_wishbone_bd_ram_n21784,
         p_wishbone_bd_ram_n21785, p_wishbone_bd_ram_n21786,
         p_wishbone_bd_ram_n21787, p_wishbone_bd_ram_n21788,
         p_wishbone_bd_ram_n21789, p_wishbone_bd_ram_n21790,
         p_wishbone_bd_ram_n21791, p_wishbone_bd_ram_n21792,
         p_wishbone_bd_ram_n21793, p_wishbone_bd_ram_n21794,
         p_wishbone_bd_ram_n21795, p_wishbone_bd_ram_n21796,
         p_wishbone_bd_ram_n21797, p_wishbone_bd_ram_n21798,
         p_wishbone_bd_ram_n21799, p_wishbone_bd_ram_n21800,
         p_wishbone_bd_ram_n21801, p_wishbone_bd_ram_n21802,
         p_wishbone_bd_ram_n21803, p_wishbone_bd_ram_n21804,
         p_wishbone_bd_ram_n21805, p_wishbone_bd_ram_n21806,
         p_wishbone_bd_ram_n21807, p_wishbone_bd_ram_n21808,
         p_wishbone_bd_ram_n21809, p_wishbone_bd_ram_n21810,
         p_wishbone_bd_ram_n21811, p_wishbone_bd_ram_n21812,
         p_wishbone_bd_ram_n21813, p_wishbone_bd_ram_n21814,
         p_wishbone_bd_ram_n21815, p_wishbone_bd_ram_n21816,
         p_wishbone_bd_ram_n21817, p_wishbone_bd_ram_n21818,
         p_wishbone_bd_ram_n21819, p_wishbone_bd_ram_n21820,
         p_wishbone_bd_ram_n21821, p_wishbone_bd_ram_n21822,
         p_wishbone_bd_ram_n21823, p_wishbone_bd_ram_n21824,
         p_wishbone_bd_ram_n21825, p_wishbone_bd_ram_n21826,
         p_wishbone_bd_ram_n21827, p_wishbone_bd_ram_n21828,
         p_wishbone_bd_ram_n21829, p_wishbone_bd_ram_n21830,
         p_wishbone_bd_ram_n21831, p_wishbone_bd_ram_n21832,
         p_wishbone_bd_ram_n21833, p_wishbone_bd_ram_n21834,
         p_wishbone_bd_ram_n21835, p_wishbone_bd_ram_n21836,
         p_wishbone_bd_ram_n21837, p_wishbone_bd_ram_n21838,
         p_wishbone_bd_ram_n21839, p_wishbone_bd_ram_n21840,
         p_wishbone_bd_ram_n21841, p_wishbone_bd_ram_n21842,
         p_wishbone_bd_ram_n21843, p_wishbone_bd_ram_n21844,
         p_wishbone_bd_ram_n21845, p_wishbone_bd_ram_n21846,
         p_wishbone_bd_ram_n21847, p_wishbone_bd_ram_n21848,
         p_wishbone_bd_ram_n21849, p_wishbone_bd_ram_n21850,
         p_wishbone_bd_ram_n21851, p_wishbone_bd_ram_n21852,
         p_wishbone_bd_ram_n21853, p_wishbone_bd_ram_n21854,
         p_wishbone_bd_ram_n21855, p_wishbone_bd_ram_n21856,
         p_wishbone_bd_ram_n21857, p_wishbone_bd_ram_n21858,
         p_wishbone_bd_ram_n21859, p_wishbone_bd_ram_n21860,
         p_wishbone_bd_ram_n21861, p_wishbone_bd_ram_n21862,
         p_wishbone_bd_ram_n21863, p_wishbone_bd_ram_n21864,
         p_wishbone_bd_ram_n21865, p_wishbone_bd_ram_n21866,
         p_wishbone_bd_ram_n21867, p_wishbone_bd_ram_n21868,
         p_wishbone_bd_ram_n21869, p_wishbone_bd_ram_n21870,
         p_wishbone_bd_ram_n21871, p_wishbone_bd_ram_n21872,
         p_wishbone_bd_ram_n21873, p_wishbone_bd_ram_n21874,
         p_wishbone_bd_ram_n21875, p_wishbone_bd_ram_n21876,
         p_wishbone_bd_ram_n21877, p_wishbone_bd_ram_n21878,
         p_wishbone_bd_ram_n21879, p_wishbone_bd_ram_n21880,
         p_wishbone_bd_ram_n21881, p_wishbone_bd_ram_n21882,
         p_wishbone_bd_ram_n21883, p_wishbone_bd_ram_n21884,
         p_wishbone_bd_ram_n21885, p_wishbone_bd_ram_n21886,
         p_wishbone_bd_ram_n21887, p_wishbone_bd_ram_n21888,
         p_wishbone_bd_ram_n21889, p_wishbone_bd_ram_n21890,
         p_wishbone_bd_ram_n21891, p_wishbone_bd_ram_n21892,
         p_wishbone_bd_ram_n21893, p_wishbone_bd_ram_n21894,
         p_wishbone_bd_ram_n21895, p_wishbone_bd_ram_n21896,
         p_wishbone_bd_ram_n21897, p_wishbone_bd_ram_n21898,
         p_wishbone_bd_ram_n21899, p_wishbone_bd_ram_n21900,
         p_wishbone_bd_ram_n21901, p_wishbone_bd_ram_n21902,
         p_wishbone_bd_ram_n21903, p_wishbone_bd_ram_n21904,
         p_wishbone_bd_ram_n21905, p_wishbone_bd_ram_n21906,
         p_wishbone_bd_ram_n21907, p_wishbone_bd_ram_n21908,
         p_wishbone_bd_ram_n21909, p_wishbone_bd_ram_n21910,
         p_wishbone_bd_ram_n21911, p_wishbone_bd_ram_n21912,
         p_wishbone_bd_ram_n21913, p_wishbone_bd_ram_n21914,
         p_wishbone_bd_ram_n21915, p_wishbone_bd_ram_n21916,
         p_wishbone_bd_ram_n21917, p_wishbone_bd_ram_n21918,
         p_wishbone_bd_ram_n21919, p_wishbone_bd_ram_n21920,
         p_wishbone_bd_ram_n21921, p_wishbone_bd_ram_n21922,
         p_wishbone_bd_ram_n21923, p_wishbone_bd_ram_n21924,
         p_wishbone_bd_ram_n21925, p_wishbone_bd_ram_n21926,
         p_wishbone_bd_ram_n21927, p_wishbone_bd_ram_n21928,
         p_wishbone_bd_ram_n21929, p_wishbone_bd_ram_n21930,
         p_wishbone_bd_ram_n21931, p_wishbone_bd_ram_n21932,
         p_wishbone_bd_ram_n21933, p_wishbone_bd_ram_n21934,
         p_wishbone_bd_ram_n21935, p_wishbone_bd_ram_n21936,
         p_wishbone_bd_ram_n21937, p_wishbone_bd_ram_n21938,
         p_wishbone_bd_ram_n21939, p_wishbone_bd_ram_n21940,
         p_wishbone_bd_ram_n21941, p_wishbone_bd_ram_n21942,
         p_wishbone_bd_ram_n21943, p_wishbone_bd_ram_n21944,
         p_wishbone_bd_ram_n21945, p_wishbone_bd_ram_n21946,
         p_wishbone_bd_ram_n21947, p_wishbone_bd_ram_n21948,
         p_wishbone_bd_ram_n21949, p_wishbone_bd_ram_n21950,
         p_wishbone_bd_ram_n21951, p_wishbone_bd_ram_n21952,
         p_wishbone_bd_ram_n21953, p_wishbone_bd_ram_n21954,
         p_wishbone_bd_ram_n21955, p_wishbone_bd_ram_n21956,
         p_wishbone_bd_ram_n21957, p_wishbone_bd_ram_n21958,
         p_wishbone_bd_ram_n21959, p_wishbone_bd_ram_n21960,
         p_wishbone_bd_ram_n21961, p_wishbone_bd_ram_n21962,
         p_wishbone_bd_ram_n21963, p_wishbone_bd_ram_n21964,
         p_wishbone_bd_ram_n21965, p_wishbone_bd_ram_n21966,
         p_wishbone_bd_ram_n21967, p_wishbone_bd_ram_n21968,
         p_wishbone_bd_ram_n21969, p_wishbone_bd_ram_n21970,
         p_wishbone_bd_ram_n21971, p_wishbone_bd_ram_n21972,
         p_wishbone_bd_ram_n21973, p_wishbone_bd_ram_n21974,
         p_wishbone_bd_ram_n21975, p_wishbone_bd_ram_n21976,
         p_wishbone_bd_ram_n21977, p_wishbone_bd_ram_n21978,
         p_wishbone_bd_ram_n21979, p_wishbone_bd_ram_n21980,
         p_wishbone_bd_ram_n21981, p_wishbone_bd_ram_n21982,
         p_wishbone_bd_ram_n21983, p_wishbone_bd_ram_n21984,
         p_wishbone_bd_ram_n21985, p_wishbone_bd_ram_n21986,
         p_wishbone_bd_ram_n21987, p_wishbone_bd_ram_n21988,
         p_wishbone_bd_ram_n21989, p_wishbone_bd_ram_n21990,
         p_wishbone_bd_ram_n21991, p_wishbone_bd_ram_n21992,
         p_wishbone_bd_ram_n21993, p_wishbone_bd_ram_n21994,
         p_wishbone_bd_ram_n21995, p_wishbone_bd_ram_n21996,
         p_wishbone_bd_ram_n21997, p_wishbone_bd_ram_n21998,
         p_wishbone_bd_ram_n21999, p_wishbone_bd_ram_n22000,
         p_wishbone_bd_ram_n22001, p_wishbone_bd_ram_n22002,
         p_wishbone_bd_ram_n22003, p_wishbone_bd_ram_n22004,
         p_wishbone_bd_ram_n22005, p_wishbone_bd_ram_n22006,
         p_wishbone_bd_ram_n22007, p_wishbone_bd_ram_n22008,
         p_wishbone_bd_ram_n22009, p_wishbone_bd_ram_n22010,
         p_wishbone_bd_ram_n22011, p_wishbone_bd_ram_n22012,
         p_wishbone_bd_ram_n22013, p_wishbone_bd_ram_n22014,
         p_wishbone_bd_ram_n22015, p_wishbone_bd_ram_n22016,
         p_wishbone_bd_ram_n22017, p_wishbone_bd_ram_n22018,
         p_wishbone_bd_ram_n22019, p_wishbone_bd_ram_n22020,
         p_wishbone_bd_ram_n22021, p_wishbone_bd_ram_n22022,
         p_wishbone_bd_ram_n22023, p_wishbone_bd_ram_n22024,
         p_wishbone_bd_ram_n22025, p_wishbone_bd_ram_n22026,
         p_wishbone_bd_ram_n22027, p_wishbone_bd_ram_n22028,
         p_wishbone_bd_ram_n22029, p_wishbone_bd_ram_n22030,
         p_wishbone_bd_ram_n22031, p_wishbone_bd_ram_n22032,
         p_wishbone_bd_ram_n22033, p_wishbone_bd_ram_n22034,
         p_wishbone_bd_ram_n22035, p_wishbone_bd_ram_n22036,
         p_wishbone_bd_ram_n22037, p_wishbone_bd_ram_n22038,
         p_wishbone_bd_ram_n22039, p_wishbone_bd_ram_n22040,
         p_wishbone_bd_ram_n22041, p_wishbone_bd_ram_n22042,
         p_wishbone_bd_ram_n22043, p_wishbone_bd_ram_n22044,
         p_wishbone_bd_ram_n22045, p_wishbone_bd_ram_n22046,
         p_wishbone_bd_ram_n22047, p_wishbone_bd_ram_n22048,
         p_wishbone_bd_ram_n22049, p_wishbone_bd_ram_n22050,
         p_wishbone_bd_ram_n22051, p_wishbone_bd_ram_n22052,
         p_wishbone_bd_ram_n22053, p_wishbone_bd_ram_n22054,
         p_wishbone_bd_ram_n22055, p_wishbone_bd_ram_n22056,
         p_wishbone_bd_ram_n22057, p_wishbone_bd_ram_n22058,
         p_wishbone_bd_ram_n22059, p_wishbone_bd_ram_n22060,
         p_wishbone_bd_ram_n22061, p_wishbone_bd_ram_n22062,
         p_wishbone_bd_ram_n22063, p_wishbone_bd_ram_n22064,
         p_wishbone_bd_ram_n22065, p_wishbone_bd_ram_n22066,
         p_wishbone_bd_ram_n22067, p_wishbone_bd_ram_n22068,
         p_wishbone_bd_ram_n22069, p_wishbone_bd_ram_n22070,
         p_wishbone_bd_ram_n22071, p_wishbone_bd_ram_n22072,
         p_wishbone_bd_ram_n22073, p_wishbone_bd_ram_n22074,
         p_wishbone_bd_ram_n22075, p_wishbone_bd_ram_n22076,
         p_wishbone_bd_ram_n22077, p_wishbone_bd_ram_n22078,
         p_wishbone_bd_ram_n22079, p_wishbone_bd_ram_n22080,
         p_wishbone_bd_ram_n22081, p_wishbone_bd_ram_n22082,
         p_wishbone_bd_ram_n22083, p_wishbone_bd_ram_n22084,
         p_wishbone_bd_ram_n22085, p_wishbone_bd_ram_n22086,
         p_wishbone_bd_ram_n22087, p_wishbone_bd_ram_n22088,
         p_wishbone_bd_ram_n22089, p_wishbone_bd_ram_n22090,
         p_wishbone_bd_ram_n22091, p_wishbone_bd_ram_n22092,
         p_wishbone_bd_ram_n22093, p_wishbone_bd_ram_n22094,
         p_wishbone_bd_ram_n22095, p_wishbone_bd_ram_n22096,
         p_wishbone_bd_ram_n22097, p_wishbone_bd_ram_n22098,
         p_wishbone_bd_ram_n22099, p_wishbone_bd_ram_n22100,
         p_wishbone_bd_ram_n22101, p_wishbone_bd_ram_n22102,
         p_wishbone_bd_ram_n22103, p_wishbone_bd_ram_n22104,
         p_wishbone_bd_ram_n22105, p_wishbone_bd_ram_n22106,
         p_wishbone_bd_ram_n22107, p_wishbone_bd_ram_n22108,
         p_wishbone_bd_ram_n22109, p_wishbone_bd_ram_n22110,
         p_wishbone_bd_ram_n22111, p_wishbone_bd_ram_n22112,
         p_wishbone_bd_ram_n22113, p_wishbone_bd_ram_n22114,
         p_wishbone_bd_ram_n22115, p_wishbone_bd_ram_n22116,
         p_wishbone_bd_ram_n22117, p_wishbone_bd_ram_n22118,
         p_wishbone_bd_ram_n22119, p_wishbone_bd_ram_n22120,
         p_wishbone_bd_ram_n22121, p_wishbone_bd_ram_n22122,
         p_wishbone_bd_ram_n22123, p_wishbone_bd_ram_n22124,
         p_wishbone_bd_ram_n22125, p_wishbone_bd_ram_n22126,
         p_wishbone_bd_ram_n22127, p_wishbone_bd_ram_n22128,
         p_wishbone_bd_ram_n22129, p_wishbone_bd_ram_n22130,
         p_wishbone_bd_ram_n22131, p_wishbone_bd_ram_n22132,
         p_wishbone_bd_ram_n22133, p_wishbone_bd_ram_n22134,
         p_wishbone_bd_ram_n22135, p_wishbone_bd_ram_n22136,
         p_wishbone_bd_ram_n22137, p_wishbone_bd_ram_n22138,
         p_wishbone_bd_ram_n22139, p_wishbone_bd_ram_n22140,
         p_wishbone_bd_ram_n22141, p_wishbone_bd_ram_n22142,
         p_wishbone_bd_ram_n22143, p_wishbone_bd_ram_n22144,
         p_wishbone_bd_ram_n22145, p_wishbone_bd_ram_n22146,
         p_wishbone_bd_ram_n22147, p_wishbone_bd_ram_n22148,
         p_wishbone_bd_ram_n22149, p_wishbone_bd_ram_n22150,
         p_wishbone_bd_ram_n22151, p_wishbone_bd_ram_n22152,
         p_wishbone_bd_ram_n22153, p_wishbone_bd_ram_n22154,
         p_wishbone_bd_ram_n22155, p_wishbone_bd_ram_n22156,
         p_wishbone_bd_ram_n22157, p_wishbone_bd_ram_n22158,
         p_wishbone_bd_ram_n22159, p_wishbone_bd_ram_n22160,
         p_wishbone_bd_ram_n22161, p_wishbone_bd_ram_n22162,
         p_wishbone_bd_ram_n22163, p_wishbone_bd_ram_n22164,
         p_wishbone_bd_ram_n22165, p_wishbone_bd_ram_n22166,
         p_wishbone_bd_ram_n22167, p_wishbone_bd_ram_n22168,
         p_wishbone_bd_ram_n22169, p_wishbone_bd_ram_n22170,
         p_wishbone_bd_ram_n22171, p_wishbone_bd_ram_n22172,
         p_wishbone_bd_ram_n22173, p_wishbone_bd_ram_n22174,
         p_wishbone_bd_ram_n22175, p_wishbone_bd_ram_n22176,
         p_wishbone_bd_ram_n22177, p_wishbone_bd_ram_n22178,
         p_wishbone_bd_ram_n22179, p_wishbone_bd_ram_n22180,
         p_wishbone_bd_ram_n22181, p_wishbone_bd_ram_n22182,
         p_wishbone_bd_ram_n22183, p_wishbone_bd_ram_n22184,
         p_wishbone_bd_ram_n22185, p_wishbone_bd_ram_n22186,
         p_wishbone_bd_ram_n22187, p_wishbone_bd_ram_n22188,
         p_wishbone_bd_ram_n22189, p_wishbone_bd_ram_n22190,
         p_wishbone_bd_ram_n22191, p_wishbone_bd_ram_n22192,
         p_wishbone_bd_ram_n22193, p_wishbone_bd_ram_n22194,
         p_wishbone_bd_ram_n22195, p_wishbone_bd_ram_n22196,
         p_wishbone_bd_ram_n22197, p_wishbone_bd_ram_n22198,
         p_wishbone_bd_ram_n22199, p_wishbone_bd_ram_n22200,
         p_wishbone_bd_ram_n22201, p_wishbone_bd_ram_n22202,
         p_wishbone_bd_ram_n22203, p_wishbone_bd_ram_n22204,
         p_wishbone_bd_ram_n22205, p_wishbone_bd_ram_n22206,
         p_wishbone_bd_ram_n22207, p_wishbone_bd_ram_n22208,
         p_wishbone_bd_ram_n22209, p_wishbone_bd_ram_n22210,
         p_wishbone_bd_ram_n22211, p_wishbone_bd_ram_n22212,
         p_wishbone_bd_ram_n22213, p_wishbone_bd_ram_n22214,
         p_wishbone_bd_ram_n22215, p_wishbone_bd_ram_n22216,
         p_wishbone_bd_ram_n22217, p_wishbone_bd_ram_n22218,
         p_wishbone_bd_ram_n22219, p_wishbone_bd_ram_n22220,
         p_wishbone_bd_ram_n22221, p_wishbone_bd_ram_n22222,
         p_wishbone_bd_ram_n22223, p_wishbone_bd_ram_n22224,
         p_wishbone_bd_ram_n22225, p_wishbone_bd_ram_n22226,
         p_wishbone_bd_ram_n22227, p_wishbone_bd_ram_n22228,
         p_wishbone_bd_ram_n22229, p_wishbone_bd_ram_n22230,
         p_wishbone_bd_ram_n22231, p_wishbone_bd_ram_n22232,
         p_wishbone_bd_ram_n22233, p_wishbone_bd_ram_n22234,
         p_wishbone_bd_ram_n22235, p_wishbone_bd_ram_n22236,
         p_wishbone_bd_ram_n22237, p_wishbone_bd_ram_n22238,
         p_wishbone_bd_ram_n22239, p_wishbone_bd_ram_n22240,
         p_wishbone_bd_ram_n22241, p_wishbone_bd_ram_n22242,
         p_wishbone_bd_ram_n22243, p_wishbone_bd_ram_n22244,
         p_wishbone_bd_ram_n22245, p_wishbone_bd_ram_n22246,
         p_wishbone_bd_ram_n22247, p_wishbone_bd_ram_n22248,
         p_wishbone_bd_ram_n22249, p_wishbone_bd_ram_n22250,
         p_wishbone_bd_ram_n22251, p_wishbone_bd_ram_n22252,
         p_wishbone_bd_ram_n22253, p_wishbone_bd_ram_n22254,
         p_wishbone_bd_ram_n22255, p_wishbone_bd_ram_n22256,
         p_wishbone_bd_ram_n22257, p_wishbone_bd_ram_n22258,
         p_wishbone_bd_ram_n22259, p_wishbone_bd_ram_n22260,
         p_wishbone_bd_ram_n22261, p_wishbone_bd_ram_n22262,
         p_wishbone_bd_ram_n22263, p_wishbone_bd_ram_n22264,
         p_wishbone_bd_ram_n22265, p_wishbone_bd_ram_n22266,
         p_wishbone_bd_ram_n22267, p_wishbone_bd_ram_n22268,
         p_wishbone_bd_ram_n22269, p_wishbone_bd_ram_n22270,
         p_wishbone_bd_ram_n22271, p_wishbone_bd_ram_n22272,
         p_wishbone_bd_ram_n22273, p_wishbone_bd_ram_n22274,
         p_wishbone_bd_ram_n22275, p_wishbone_bd_ram_n22276,
         p_wishbone_bd_ram_n22277, p_wishbone_bd_ram_n22278,
         p_wishbone_bd_ram_n22279, p_wishbone_bd_ram_n22280,
         p_wishbone_bd_ram_n22281, p_wishbone_bd_ram_n22282,
         p_wishbone_bd_ram_n22283, p_wishbone_bd_ram_n22284,
         p_wishbone_bd_ram_n22285, p_wishbone_bd_ram_n22286,
         p_wishbone_bd_ram_n22287, p_wishbone_bd_ram_n22288,
         p_wishbone_bd_ram_n22289, p_wishbone_bd_ram_n22290,
         p_wishbone_bd_ram_n22291, p_wishbone_bd_ram_n22292,
         p_wishbone_bd_ram_n22293, p_wishbone_bd_ram_n22294,
         p_wishbone_bd_ram_n22295, p_wishbone_bd_ram_n22296,
         p_wishbone_bd_ram_n22297, p_wishbone_bd_ram_n22298,
         p_wishbone_bd_ram_n22299, p_wishbone_bd_ram_n22300,
         p_wishbone_bd_ram_n22301, p_wishbone_bd_ram_n22302,
         p_wishbone_bd_ram_n22303, p_wishbone_bd_ram_n22304,
         p_wishbone_bd_ram_n22305, p_wishbone_bd_ram_n22306,
         p_wishbone_bd_ram_n22307, p_wishbone_bd_ram_n22308,
         p_wishbone_bd_ram_n22309, p_wishbone_bd_ram_n22310,
         p_wishbone_bd_ram_n22311, p_wishbone_bd_ram_n22312,
         p_wishbone_bd_ram_n22313, p_wishbone_bd_ram_n22314,
         p_wishbone_bd_ram_n22315, p_wishbone_bd_ram_n22316,
         p_wishbone_bd_ram_n22317, p_wishbone_bd_ram_n22318,
         p_wishbone_bd_ram_n22319, p_wishbone_bd_ram_n22320,
         p_wishbone_bd_ram_n22321, p_wishbone_bd_ram_n22322,
         p_wishbone_bd_ram_n22323, p_wishbone_bd_ram_n22324,
         p_wishbone_bd_ram_n22325, p_wishbone_bd_ram_n22326,
         p_wishbone_bd_ram_n22327, p_wishbone_bd_ram_n22328,
         p_wishbone_bd_ram_n22329, p_wishbone_bd_ram_n22330,
         p_wishbone_bd_ram_n22331, p_wishbone_bd_ram_n22332,
         p_wishbone_bd_ram_n22333, p_wishbone_bd_ram_n22334,
         p_wishbone_bd_ram_n22335, p_wishbone_bd_ram_n22336,
         p_wishbone_bd_ram_n22337, p_wishbone_bd_ram_n22338,
         p_wishbone_bd_ram_n22339, p_wishbone_bd_ram_n22340,
         p_wishbone_bd_ram_n22341, p_wishbone_bd_ram_n22342,
         p_wishbone_bd_ram_n22343, p_wishbone_bd_ram_n22344,
         p_wishbone_bd_ram_n22345, p_wishbone_bd_ram_n22346,
         p_wishbone_bd_ram_n22347, p_wishbone_bd_ram_n22348,
         p_wishbone_bd_ram_n22349, p_wishbone_bd_ram_n22350,
         p_wishbone_bd_ram_n22351, p_wishbone_bd_ram_n22352,
         p_wishbone_bd_ram_n22353, p_wishbone_bd_ram_n22354,
         p_wishbone_bd_ram_n22355, p_wishbone_bd_ram_n22356,
         p_wishbone_bd_ram_n22357, p_wishbone_bd_ram_n22358,
         p_wishbone_bd_ram_n22359, p_wishbone_bd_ram_n22360,
         p_wishbone_bd_ram_n22361, p_wishbone_bd_ram_n22362,
         p_wishbone_bd_ram_n22363, p_wishbone_bd_ram_n22364,
         p_wishbone_bd_ram_n22365, p_wishbone_bd_ram_n22366,
         p_wishbone_bd_ram_n22367, p_wishbone_bd_ram_n22368,
         p_wishbone_bd_ram_n22369, p_wishbone_bd_ram_n22370,
         p_wishbone_bd_ram_n22371, p_wishbone_bd_ram_n22372,
         p_wishbone_bd_ram_n22373, p_wishbone_bd_ram_n22374,
         p_wishbone_bd_ram_n22375, p_wishbone_bd_ram_n22376,
         p_wishbone_bd_ram_n22377, p_wishbone_bd_ram_n22378,
         p_wishbone_bd_ram_n22379, p_wishbone_bd_ram_n22380,
         p_wishbone_bd_ram_n22381, p_wishbone_bd_ram_n22382,
         p_wishbone_bd_ram_n22383, p_wishbone_bd_ram_n22384,
         p_wishbone_bd_ram_n22385, p_wishbone_bd_ram_n22386,
         p_wishbone_bd_ram_n22387, p_wishbone_bd_ram_n22388,
         p_wishbone_bd_ram_n22389, p_wishbone_bd_ram_n22390,
         p_wishbone_bd_ram_n22391, p_wishbone_bd_ram_n22392,
         p_wishbone_bd_ram_n22393, p_wishbone_bd_ram_n22394,
         p_wishbone_bd_ram_n22395, p_wishbone_bd_ram_n22396,
         p_wishbone_bd_ram_n22397, p_wishbone_bd_ram_n22398,
         p_wishbone_bd_ram_n22399, p_wishbone_bd_ram_n22400,
         p_wishbone_bd_ram_n22401, p_wishbone_bd_ram_n22402,
         p_wishbone_bd_ram_n22403, p_wishbone_bd_ram_n22404,
         p_wishbone_bd_ram_n22405, p_wishbone_bd_ram_n22406,
         p_wishbone_bd_ram_n22407, p_wishbone_bd_ram_n22408,
         p_wishbone_bd_ram_n22409, p_wishbone_bd_ram_n22410,
         p_wishbone_bd_ram_n22411, p_wishbone_bd_ram_n22412,
         p_wishbone_bd_ram_n22413, p_wishbone_bd_ram_n22414,
         p_wishbone_bd_ram_n22415, p_wishbone_bd_ram_n22416,
         p_wishbone_bd_ram_n22417, p_wishbone_bd_ram_n22418,
         p_wishbone_bd_ram_n22419, p_wishbone_bd_ram_n22420,
         p_wishbone_bd_ram_n22421, p_wishbone_bd_ram_n22422,
         p_wishbone_bd_ram_n22423, p_wishbone_bd_ram_n22424,
         p_wishbone_bd_ram_n22425, p_wishbone_bd_ram_n22426,
         p_wishbone_bd_ram_n22427, p_wishbone_bd_ram_n22428,
         p_wishbone_bd_ram_n22429, p_wishbone_bd_ram_n22430,
         p_wishbone_bd_ram_n22431, p_wishbone_bd_ram_n22432,
         p_wishbone_bd_ram_n22433, p_wishbone_bd_ram_n22434,
         p_wishbone_bd_ram_n22435, p_wishbone_bd_ram_n22436,
         p_wishbone_bd_ram_n22437, p_wishbone_bd_ram_n22438,
         p_wishbone_bd_ram_n22439, p_wishbone_bd_ram_n22440,
         p_wishbone_bd_ram_n22441, p_wishbone_bd_ram_n22442,
         p_wishbone_bd_ram_n22443, p_wishbone_bd_ram_n22444,
         p_wishbone_bd_ram_n22445, p_wishbone_bd_ram_n22446,
         p_wishbone_bd_ram_n22447, p_wishbone_bd_ram_n22448,
         p_wishbone_bd_ram_n22449, p_wishbone_bd_ram_n22450,
         p_wishbone_bd_ram_n22451, p_wishbone_bd_ram_n22452,
         p_wishbone_bd_ram_n22453, p_wishbone_bd_ram_n22454,
         p_wishbone_bd_ram_n22455, p_wishbone_bd_ram_n22456,
         p_wishbone_bd_ram_n22457, p_wishbone_bd_ram_n22458,
         p_wishbone_bd_ram_n22459, p_wishbone_bd_ram_n22460,
         p_wishbone_bd_ram_n22461, p_wishbone_bd_ram_n22462,
         p_wishbone_bd_ram_n22463, p_wishbone_bd_ram_n22464,
         p_wishbone_bd_ram_n22465, p_wishbone_bd_ram_n22466,
         p_wishbone_bd_ram_n22467, p_wishbone_bd_ram_n22468,
         p_wishbone_bd_ram_n22469, p_wishbone_bd_ram_n22470,
         p_wishbone_bd_ram_n22471, p_wishbone_bd_ram_n22472,
         p_wishbone_bd_ram_n22473, p_wishbone_bd_ram_n22474,
         p_wishbone_bd_ram_n22475, p_wishbone_bd_ram_n22476,
         p_wishbone_bd_ram_n22477, p_wishbone_bd_ram_n22478,
         p_wishbone_bd_ram_n22479, p_wishbone_bd_ram_n22480,
         p_wishbone_bd_ram_n22481, p_wishbone_bd_ram_n22482,
         p_wishbone_bd_ram_n22483, p_wishbone_bd_ram_n22484,
         p_wishbone_bd_ram_n22485, p_wishbone_bd_ram_n22486,
         p_wishbone_bd_ram_n22487, p_wishbone_bd_ram_n22488,
         p_wishbone_bd_ram_n22489, p_wishbone_bd_ram_n22490,
         p_wishbone_bd_ram_n22491, p_wishbone_bd_ram_n22492,
         p_wishbone_bd_ram_n22493, p_wishbone_bd_ram_n22494,
         p_wishbone_bd_ram_n22495, p_wishbone_bd_ram_n22496,
         p_wishbone_bd_ram_n22497, p_wishbone_bd_ram_n22498,
         p_wishbone_bd_ram_n22499, p_wishbone_bd_ram_n22500,
         p_wishbone_bd_ram_n22501, p_wishbone_bd_ram_n22502,
         p_wishbone_bd_ram_n22503, p_wishbone_bd_ram_n22504,
         p_wishbone_bd_ram_n22505, p_wishbone_bd_ram_n22506,
         p_wishbone_bd_ram_n22507, p_wishbone_bd_ram_n22508,
         p_wishbone_bd_ram_n22509, p_wishbone_bd_ram_n22510,
         p_wishbone_bd_ram_n22511, p_wishbone_bd_ram_n22512,
         p_wishbone_bd_ram_n22513, p_wishbone_bd_ram_n22514,
         p_wishbone_bd_ram_n22515, p_wishbone_bd_ram_n22516,
         p_wishbone_bd_ram_n22517, p_wishbone_bd_ram_n22518,
         p_wishbone_bd_ram_n22519, p_wishbone_bd_ram_n22520,
         p_wishbone_bd_ram_n22521, p_wishbone_bd_ram_n22522,
         p_wishbone_bd_ram_n22523, p_wishbone_bd_ram_n22524,
         p_wishbone_bd_ram_n22525, p_wishbone_bd_ram_n22526,
         p_wishbone_bd_ram_n22527, p_wishbone_bd_ram_n22528,
         p_wishbone_bd_ram_n22529, p_wishbone_bd_ram_n22530,
         p_wishbone_bd_ram_n22531, p_wishbone_bd_ram_n22532,
         p_wishbone_bd_ram_n22533, p_wishbone_bd_ram_n22534,
         p_wishbone_bd_ram_n22535, p_wishbone_bd_ram_n22536,
         p_wishbone_bd_ram_n22537, p_wishbone_bd_ram_n22538,
         p_wishbone_bd_ram_n22539, p_wishbone_bd_ram_n22540,
         p_wishbone_bd_ram_n22541, p_wishbone_bd_ram_n22542,
         p_wishbone_bd_ram_n22543, p_wishbone_bd_ram_n22544,
         p_wishbone_bd_ram_n22545, p_wishbone_bd_ram_n22546,
         p_wishbone_bd_ram_n22547, p_wishbone_bd_ram_n22548,
         p_wishbone_bd_ram_n22549, p_wishbone_bd_ram_n22550,
         p_wishbone_bd_ram_n22551, p_wishbone_bd_ram_n22552,
         p_wishbone_bd_ram_n22553, p_wishbone_bd_ram_n22554,
         p_wishbone_bd_ram_n22555, p_wishbone_bd_ram_n22556,
         p_wishbone_bd_ram_n22557, p_wishbone_bd_ram_n22558,
         p_wishbone_bd_ram_n22559, p_wishbone_bd_ram_n22560,
         p_wishbone_bd_ram_n22561, p_wishbone_bd_ram_n22562,
         p_wishbone_bd_ram_n22563, p_wishbone_bd_ram_n22564,
         p_wishbone_bd_ram_n22565, p_wishbone_bd_ram_n22566,
         p_wishbone_bd_ram_n22567, p_wishbone_bd_ram_n22568,
         p_wishbone_bd_ram_n22569, p_wishbone_bd_ram_n22570,
         p_wishbone_bd_ram_n22571, p_wishbone_bd_ram_n22572,
         p_wishbone_bd_ram_n22573, p_wishbone_bd_ram_n22574,
         p_wishbone_bd_ram_n22575, p_wishbone_bd_ram_n22576,
         p_wishbone_bd_ram_n22577, p_wishbone_bd_ram_n22578,
         p_wishbone_bd_ram_n22579, p_wishbone_bd_ram_n22580,
         p_wishbone_bd_ram_n22581, p_wishbone_bd_ram_n22582,
         p_wishbone_bd_ram_n22583, p_wishbone_bd_ram_n22584,
         p_wishbone_bd_ram_n22585, p_wishbone_bd_ram_n22586,
         p_wishbone_bd_ram_n22587, p_wishbone_bd_ram_n22588,
         p_wishbone_bd_ram_n22589, p_wishbone_bd_ram_n22590,
         p_wishbone_bd_ram_n22591, p_wishbone_bd_ram_n22592,
         p_wishbone_bd_ram_n22593, p_wishbone_bd_ram_n22594,
         p_wishbone_bd_ram_n22595, p_wishbone_bd_ram_n22596,
         p_wishbone_bd_ram_n22597, p_wishbone_bd_ram_n22598,
         p_wishbone_bd_ram_n22599, p_wishbone_bd_ram_n22600,
         p_wishbone_bd_ram_n22601, p_wishbone_bd_ram_n22602,
         p_wishbone_bd_ram_n22603, p_wishbone_bd_ram_n22604,
         p_wishbone_bd_ram_n22605, p_wishbone_bd_ram_n22606,
         p_wishbone_bd_ram_n22607, p_wishbone_bd_ram_n22608,
         p_wishbone_bd_ram_n22609, p_wishbone_bd_ram_n22610,
         p_wishbone_bd_ram_n22611, p_wishbone_bd_ram_n22612,
         p_wishbone_bd_ram_n22613, p_wishbone_bd_ram_n22614,
         p_wishbone_bd_ram_n22615, p_wishbone_bd_ram_n22616,
         p_wishbone_bd_ram_n22617, p_wishbone_bd_ram_n22618,
         p_wishbone_bd_ram_n22619, p_wishbone_bd_ram_n22620,
         p_wishbone_bd_ram_n22621, p_wishbone_bd_ram_n22622,
         p_wishbone_bd_ram_n22623, p_wishbone_bd_ram_n22624,
         p_wishbone_bd_ram_n22625, p_wishbone_bd_ram_n22626,
         p_wishbone_bd_ram_n22627, p_wishbone_bd_ram_n22628,
         p_wishbone_bd_ram_n22629, p_wishbone_bd_ram_n22630,
         p_wishbone_bd_ram_n22631, p_wishbone_bd_ram_n22632,
         p_wishbone_bd_ram_n22633, p_wishbone_bd_ram_n22634,
         p_wishbone_bd_ram_n22635, p_wishbone_bd_ram_n22636,
         p_wishbone_bd_ram_n22637, p_wishbone_bd_ram_n22638,
         p_wishbone_bd_ram_n22639, p_wishbone_bd_ram_n22640,
         p_wishbone_bd_ram_n22641, p_wishbone_bd_ram_n22642,
         p_wishbone_bd_ram_n22643, p_wishbone_bd_ram_n22644,
         p_wishbone_bd_ram_n22645, p_wishbone_bd_ram_n22646,
         p_wishbone_bd_ram_n22647, p_wishbone_bd_ram_n22648,
         p_wishbone_bd_ram_n22649, p_wishbone_bd_ram_n22650,
         p_wishbone_bd_ram_n22651, p_wishbone_bd_ram_n22652,
         p_wishbone_bd_ram_n22653, p_wishbone_bd_ram_n22654,
         p_wishbone_bd_ram_n22655, p_wishbone_bd_ram_n22656,
         p_wishbone_bd_ram_n22657, p_wishbone_bd_ram_n22658,
         p_wishbone_bd_ram_n22659, p_wishbone_bd_ram_n22660,
         p_wishbone_bd_ram_n22661, p_wishbone_bd_ram_n22662,
         p_wishbone_bd_ram_n22663, p_wishbone_bd_ram_n22664,
         p_wishbone_bd_ram_n22665, p_wishbone_bd_ram_n22666,
         p_wishbone_bd_ram_n22667, p_wishbone_bd_ram_n22668,
         p_wishbone_bd_ram_n22669, p_wishbone_bd_ram_n22670,
         p_wishbone_bd_ram_n22671, p_wishbone_bd_ram_n22672,
         p_wishbone_bd_ram_n22673, p_wishbone_bd_ram_n22674,
         p_wishbone_bd_ram_n22675, p_wishbone_bd_ram_n22676,
         p_wishbone_bd_ram_n22677, p_wishbone_bd_ram_n22678,
         p_wishbone_bd_ram_n22679, p_wishbone_bd_ram_n22680,
         p_wishbone_bd_ram_n22681, p_wishbone_bd_ram_n22682,
         p_wishbone_bd_ram_n22683, p_wishbone_bd_ram_n22684,
         p_wishbone_bd_ram_n22685, p_wishbone_bd_ram_n22686,
         p_wishbone_bd_ram_n22687, p_wishbone_bd_ram_n22688,
         p_wishbone_bd_ram_n22689, p_wishbone_bd_ram_n22690,
         p_wishbone_bd_ram_n22691, p_wishbone_bd_ram_n22692,
         p_wishbone_bd_ram_n22693, p_wishbone_bd_ram_n22694,
         p_wishbone_bd_ram_n22695, p_wishbone_bd_ram_n22696,
         p_wishbone_bd_ram_n22697, p_wishbone_bd_ram_n22698,
         p_wishbone_bd_ram_n22699, p_wishbone_bd_ram_n22700,
         p_wishbone_bd_ram_n22701, p_wishbone_bd_ram_n22702,
         p_wishbone_bd_ram_n22703, p_wishbone_bd_ram_n22704,
         p_wishbone_bd_ram_n22705, p_wishbone_bd_ram_n22706,
         p_wishbone_bd_ram_n22707, p_wishbone_bd_ram_n22708,
         p_wishbone_bd_ram_n22709, p_wishbone_bd_ram_n22710,
         p_wishbone_bd_ram_n22711, p_wishbone_bd_ram_n22712,
         p_wishbone_bd_ram_n22713, p_wishbone_bd_ram_n22714,
         p_wishbone_bd_ram_n22715, p_wishbone_bd_ram_n22716,
         p_wishbone_bd_ram_n22717, p_wishbone_bd_ram_n22718,
         p_wishbone_bd_ram_n22719, p_wishbone_bd_ram_n22720,
         p_wishbone_bd_ram_n22721, p_wishbone_bd_ram_n22722,
         p_wishbone_bd_ram_n22723, p_wishbone_bd_ram_n22724,
         p_wishbone_bd_ram_n22725, p_wishbone_bd_ram_n22726,
         p_wishbone_bd_ram_n22727, p_wishbone_bd_ram_n22728,
         p_wishbone_bd_ram_n22729, p_wishbone_bd_ram_n22730,
         p_wishbone_bd_ram_n22731, p_wishbone_bd_ram_n22732,
         p_wishbone_bd_ram_n22733, p_wishbone_bd_ram_n22734,
         p_wishbone_bd_ram_n22735, p_wishbone_bd_ram_n22736,
         p_wishbone_bd_ram_n22737, p_wishbone_bd_ram_n22738,
         p_wishbone_bd_ram_n22739, p_wishbone_bd_ram_n22740,
         p_wishbone_bd_ram_n22741, p_wishbone_bd_ram_n22742,
         p_wishbone_bd_ram_n22743, p_wishbone_bd_ram_n22744,
         p_wishbone_bd_ram_n22745, p_wishbone_bd_ram_n22746,
         p_wishbone_bd_ram_n22747, p_wishbone_bd_ram_n22748,
         p_wishbone_bd_ram_n22749, p_wishbone_bd_ram_n22750,
         p_wishbone_bd_ram_n22751, p_wishbone_bd_ram_n22752,
         p_wishbone_bd_ram_n22753, p_wishbone_bd_ram_n22754,
         p_wishbone_bd_ram_n22755, p_wishbone_bd_ram_n22756,
         p_wishbone_bd_ram_n22757, p_wishbone_bd_ram_n22758,
         p_wishbone_bd_ram_n22759, p_wishbone_bd_ram_n22760,
         p_wishbone_bd_ram_n22761, p_wishbone_bd_ram_n22762,
         p_wishbone_bd_ram_n22763, p_wishbone_bd_ram_n22764,
         p_wishbone_bd_ram_n22765, p_wishbone_bd_ram_n22766,
         p_wishbone_bd_ram_n22767, p_wishbone_bd_ram_n22768,
         p_wishbone_bd_ram_n22769, p_wishbone_bd_ram_n22770,
         p_wishbone_bd_ram_n22771, p_wishbone_bd_ram_n22772,
         p_wishbone_bd_ram_n22773, p_wishbone_bd_ram_n22774,
         p_wishbone_bd_ram_n22775, p_wishbone_bd_ram_n22776,
         p_wishbone_bd_ram_n22777, p_wishbone_bd_ram_n22778,
         p_wishbone_bd_ram_n22779, p_wishbone_bd_ram_n22780,
         p_wishbone_bd_ram_n22781, p_wishbone_bd_ram_n22782,
         p_wishbone_bd_ram_n22783, p_wishbone_bd_ram_n22784,
         p_wishbone_bd_ram_n22785, p_wishbone_bd_ram_n22786,
         p_wishbone_bd_ram_n22787, p_wishbone_bd_ram_n22788,
         p_wishbone_bd_ram_n22789, p_wishbone_bd_ram_n22790,
         p_wishbone_bd_ram_n22791, p_wishbone_bd_ram_n22792,
         p_wishbone_bd_ram_n22793, p_wishbone_bd_ram_n22794,
         p_wishbone_bd_ram_n22795, p_wishbone_bd_ram_n22796,
         p_wishbone_bd_ram_n22797, p_wishbone_bd_ram_n22798,
         p_wishbone_bd_ram_n22799, p_wishbone_bd_ram_n22800,
         p_wishbone_bd_ram_n22801, p_wishbone_bd_ram_n22802,
         p_wishbone_bd_ram_n22803, p_wishbone_bd_ram_n22804,
         p_wishbone_bd_ram_n22805, p_wishbone_bd_ram_n22806,
         p_wishbone_bd_ram_n22807, p_wishbone_bd_ram_n22808,
         p_wishbone_bd_ram_n22809, p_wishbone_bd_ram_n22810,
         p_wishbone_bd_ram_n22811, p_wishbone_bd_ram_n22812,
         p_wishbone_bd_ram_n22813, p_wishbone_bd_ram_n22814,
         p_wishbone_bd_ram_n22815, p_wishbone_bd_ram_n22816,
         p_wishbone_bd_ram_n22817, p_wishbone_bd_ram_n22818,
         p_wishbone_bd_ram_n22819, p_wishbone_bd_ram_n22820,
         p_wishbone_bd_ram_n22821, p_wishbone_bd_ram_n22822,
         p_wishbone_bd_ram_n22823, p_wishbone_bd_ram_n22824,
         p_wishbone_bd_ram_n22825, p_wishbone_bd_ram_n22826,
         p_wishbone_bd_ram_n22827, p_wishbone_bd_ram_n22828,
         p_wishbone_bd_ram_n22829, p_wishbone_bd_ram_n22830,
         p_wishbone_bd_ram_n22831, p_wishbone_bd_ram_n22832,
         p_wishbone_bd_ram_n22833, p_wishbone_bd_ram_n22834,
         p_wishbone_bd_ram_n22835, p_wishbone_bd_ram_n22836,
         p_wishbone_bd_ram_n22837, p_wishbone_bd_ram_n22838,
         p_wishbone_bd_ram_n22839, p_wishbone_bd_ram_n22840,
         p_wishbone_bd_ram_n22841, p_wishbone_bd_ram_n22842,
         p_wishbone_bd_ram_n22843, p_wishbone_bd_ram_n22844,
         p_wishbone_bd_ram_n22845, p_wishbone_bd_ram_n22846,
         p_wishbone_bd_ram_n22847, p_wishbone_bd_ram_n22848,
         p_wishbone_bd_ram_n22849, p_wishbone_bd_ram_n22850,
         p_wishbone_bd_ram_n22851, p_wishbone_bd_ram_n22852,
         p_wishbone_bd_ram_n22853, p_wishbone_bd_ram_n22854,
         p_wishbone_bd_ram_n22855, p_wishbone_bd_ram_n22856,
         p_wishbone_bd_ram_n22857, p_wishbone_bd_ram_n22858,
         p_wishbone_bd_ram_n22859, p_wishbone_bd_ram_n22860,
         p_wishbone_bd_ram_n22861, p_wishbone_bd_ram_n22862,
         p_wishbone_bd_ram_n22863, p_wishbone_bd_ram_n22864,
         p_wishbone_bd_ram_n22865, p_wishbone_bd_ram_n22866,
         p_wishbone_bd_ram_n22867, p_wishbone_bd_ram_n22868,
         p_wishbone_bd_ram_n22869, p_wishbone_bd_ram_n22870,
         p_wishbone_bd_ram_n22871, p_wishbone_bd_ram_n22872,
         p_wishbone_bd_ram_n22873, p_wishbone_bd_ram_n22874,
         p_wishbone_bd_ram_n22875, p_wishbone_bd_ram_n22876,
         p_wishbone_bd_ram_n22877, p_wishbone_bd_ram_n22878,
         p_wishbone_bd_ram_n22879, p_wishbone_bd_ram_n22880,
         p_wishbone_bd_ram_n22881, p_wishbone_bd_ram_n22882,
         p_wishbone_bd_ram_n22883, p_wishbone_bd_ram_n22884,
         p_wishbone_bd_ram_n22885, p_wishbone_bd_ram_n22886,
         p_wishbone_bd_ram_n22887, p_wishbone_bd_ram_n22888,
         p_wishbone_bd_ram_n22889, p_wishbone_bd_ram_n22890,
         p_wishbone_bd_ram_n22891, p_wishbone_bd_ram_n22892,
         p_wishbone_bd_ram_n22893, p_wishbone_bd_ram_n22894,
         p_wishbone_bd_ram_n22895, p_wishbone_bd_ram_n22896,
         p_wishbone_bd_ram_n22897, p_wishbone_bd_ram_n22898,
         p_wishbone_bd_ram_n22899, p_wishbone_bd_ram_n22900,
         p_wishbone_bd_ram_n22901, p_wishbone_bd_ram_n22902,
         p_wishbone_bd_ram_n22903, p_wishbone_bd_ram_n22904,
         p_wishbone_bd_ram_n22905, p_wishbone_bd_ram_n22906,
         p_wishbone_bd_ram_n22907, p_wishbone_bd_ram_n22908,
         p_wishbone_bd_ram_n22909, p_wishbone_bd_ram_n22910,
         p_wishbone_bd_ram_n22911, p_wishbone_bd_ram_n22912,
         p_wishbone_bd_ram_n22913, p_wishbone_bd_ram_n22914,
         p_wishbone_bd_ram_n22915, p_wishbone_bd_ram_n22916,
         p_wishbone_bd_ram_n22917, p_wishbone_bd_ram_n22918,
         p_wishbone_bd_ram_n22919, p_wishbone_bd_ram_n22920,
         p_wishbone_bd_ram_n22921, p_wishbone_bd_ram_n22922,
         p_wishbone_bd_ram_n22923, p_wishbone_bd_ram_n22924,
         p_wishbone_bd_ram_n22925, p_wishbone_bd_ram_n22926,
         p_wishbone_bd_ram_n22927, p_wishbone_bd_ram_n22928,
         p_wishbone_bd_ram_n22929, p_wishbone_bd_ram_n22930,
         p_wishbone_bd_ram_n22931, p_wishbone_bd_ram_n22932,
         p_wishbone_bd_ram_n22933, p_wishbone_bd_ram_n22934,
         p_wishbone_bd_ram_n22935, p_wishbone_bd_ram_n22936,
         p_wishbone_bd_ram_n22937, p_wishbone_bd_ram_n22938,
         p_wishbone_bd_ram_n22939, p_wishbone_bd_ram_n22940,
         p_wishbone_bd_ram_n22941, p_wishbone_bd_ram_n22942,
         p_wishbone_bd_ram_n22943, p_wishbone_bd_ram_n22944,
         p_wishbone_bd_ram_n22945, p_wishbone_bd_ram_n22946,
         p_wishbone_bd_ram_n22947, p_wishbone_bd_ram_n22948,
         p_wishbone_bd_ram_n22949, p_wishbone_bd_ram_n22950,
         p_wishbone_bd_ram_n22951, p_wishbone_bd_ram_n22952,
         p_wishbone_bd_ram_n22953, p_wishbone_bd_ram_n22954,
         p_wishbone_bd_ram_n22955, p_wishbone_bd_ram_n22956,
         p_wishbone_bd_ram_n22957, p_wishbone_bd_ram_n22958,
         p_wishbone_bd_ram_n22959, p_wishbone_bd_ram_n22960,
         p_wishbone_bd_ram_n22961, p_wishbone_bd_ram_n22962,
         p_wishbone_bd_ram_n22963, p_wishbone_bd_ram_n22964,
         p_wishbone_bd_ram_n22965, p_wishbone_bd_ram_n22966,
         p_wishbone_bd_ram_n22967, p_wishbone_bd_ram_n22968,
         p_wishbone_bd_ram_n22969, p_wishbone_bd_ram_n22970,
         p_wishbone_bd_ram_n22971, p_wishbone_bd_ram_n22972,
         p_wishbone_bd_ram_n22973, p_wishbone_bd_ram_n22974,
         p_wishbone_bd_ram_n22975, p_wishbone_bd_ram_n22976,
         p_wishbone_bd_ram_n22977, p_wishbone_bd_ram_n22978,
         p_wishbone_bd_ram_n22979, p_wishbone_bd_ram_n22980,
         p_wishbone_bd_ram_n22981, p_wishbone_bd_ram_n22982,
         p_wishbone_bd_ram_n22983, p_wishbone_bd_ram_n22984,
         p_wishbone_bd_ram_n22985, p_wishbone_bd_ram_n22986,
         p_wishbone_bd_ram_n22987, p_wishbone_bd_ram_n22988,
         p_wishbone_bd_ram_n22989, p_wishbone_bd_ram_n22990,
         p_wishbone_bd_ram_n22991, p_wishbone_bd_ram_n22992,
         p_wishbone_bd_ram_n22993, p_wishbone_bd_ram_n22994,
         p_wishbone_bd_ram_n22995, p_wishbone_bd_ram_n22996,
         p_wishbone_bd_ram_n22997, p_wishbone_bd_ram_n22998,
         p_wishbone_bd_ram_n22999, p_wishbone_bd_ram_n23000,
         p_wishbone_bd_ram_n23001, p_wishbone_bd_ram_n23002,
         p_wishbone_bd_ram_n23003, p_wishbone_bd_ram_n23004,
         p_wishbone_bd_ram_n23005, p_wishbone_bd_ram_n23006,
         p_wishbone_bd_ram_n23007, p_wishbone_bd_ram_n23008,
         p_wishbone_bd_ram_n23009, p_wishbone_bd_ram_n23010,
         p_wishbone_bd_ram_n23011, p_wishbone_bd_ram_n23012,
         p_wishbone_bd_ram_n23013, p_wishbone_bd_ram_n23014,
         p_wishbone_bd_ram_n23015, p_wishbone_bd_ram_n23016,
         p_wishbone_bd_ram_n23017, p_wishbone_bd_ram_n23018,
         p_wishbone_bd_ram_n23019, p_wishbone_bd_ram_n23020,
         p_wishbone_bd_ram_n23021, p_wishbone_bd_ram_n23022,
         p_wishbone_bd_ram_n23023, p_wishbone_bd_ram_n23024,
         p_wishbone_bd_ram_n23025, p_wishbone_bd_ram_n23026,
         p_wishbone_bd_ram_n23027, p_wishbone_bd_ram_n23028,
         p_wishbone_bd_ram_n23029, p_wishbone_bd_ram_n23030,
         p_wishbone_bd_ram_n23031, p_wishbone_bd_ram_n23032,
         p_wishbone_bd_ram_n23033, p_wishbone_bd_ram_n23034,
         p_wishbone_bd_ram_n23035, p_wishbone_bd_ram_n23036,
         p_wishbone_bd_ram_n23037, p_wishbone_bd_ram_n23038,
         p_wishbone_bd_ram_n23039, p_wishbone_bd_ram_n23040,
         p_wishbone_bd_ram_n23041, p_wishbone_bd_ram_n23042,
         p_wishbone_bd_ram_n23043, p_wishbone_bd_ram_n23044,
         p_wishbone_bd_ram_n23045, p_wishbone_bd_ram_n23046,
         p_wishbone_bd_ram_n23047, p_wishbone_bd_ram_n23048,
         p_wishbone_bd_ram_n23049, p_wishbone_bd_ram_n23050,
         p_wishbone_bd_ram_n23051, p_wishbone_bd_ram_n23052,
         p_wishbone_bd_ram_n23053, p_wishbone_bd_ram_n23054,
         p_wishbone_bd_ram_n23055, p_wishbone_bd_ram_n23056,
         p_wishbone_bd_ram_n23057, p_wishbone_bd_ram_n23058,
         p_wishbone_bd_ram_n23059, p_wishbone_bd_ram_n23060,
         p_wishbone_bd_ram_n23061, p_wishbone_bd_ram_n23062,
         p_wishbone_bd_ram_n23063, p_wishbone_bd_ram_n23064,
         p_wishbone_bd_ram_n23065, p_wishbone_bd_ram_n23066,
         p_wishbone_bd_ram_n23067, p_wishbone_bd_ram_n23068,
         p_wishbone_bd_ram_n23069, p_wishbone_bd_ram_n23070,
         p_wishbone_bd_ram_n23071, p_wishbone_bd_ram_n23072,
         p_wishbone_bd_ram_n23073, p_wishbone_bd_ram_n23074,
         p_wishbone_bd_ram_n23075, p_wishbone_bd_ram_n23076,
         p_wishbone_bd_ram_n23077, p_wishbone_bd_ram_n23078,
         p_wishbone_bd_ram_n23079, p_wishbone_bd_ram_n23080,
         p_wishbone_bd_ram_n23081, p_wishbone_bd_ram_n23082,
         p_wishbone_bd_ram_n23083, p_wishbone_bd_ram_n23084,
         p_wishbone_bd_ram_n23085, p_wishbone_bd_ram_n23086,
         p_wishbone_bd_ram_n23087, p_wishbone_bd_ram_n23088,
         p_wishbone_bd_ram_n23089, p_wishbone_bd_ram_n23090,
         p_wishbone_bd_ram_n23091, p_wishbone_bd_ram_n23092,
         p_wishbone_bd_ram_n23093, p_wishbone_bd_ram_n23094,
         p_wishbone_bd_ram_n23095, p_wishbone_bd_ram_n23096,
         p_wishbone_bd_ram_n23097, p_wishbone_bd_ram_n23098,
         p_wishbone_bd_ram_n23099, p_wishbone_bd_ram_n23100,
         p_wishbone_bd_ram_n23101, p_wishbone_bd_ram_n23102,
         p_wishbone_bd_ram_n23103, p_wishbone_bd_ram_n23104,
         p_wishbone_bd_ram_n23105, p_wishbone_bd_ram_n23106,
         p_wishbone_bd_ram_n23107, p_wishbone_bd_ram_n23108,
         p_wishbone_bd_ram_n23109, p_wishbone_bd_ram_n23110,
         p_wishbone_bd_ram_n23111, p_wishbone_bd_ram_n23112,
         p_wishbone_bd_ram_n23113, p_wishbone_bd_ram_n23114,
         p_wishbone_bd_ram_n23115, p_wishbone_bd_ram_n23116,
         p_wishbone_bd_ram_n23117, p_wishbone_bd_ram_n23118,
         p_wishbone_bd_ram_n23119, p_wishbone_bd_ram_n23120,
         p_wishbone_bd_ram_n23121, p_wishbone_bd_ram_n23122,
         p_wishbone_bd_ram_n23123, p_wishbone_bd_ram_n23124,
         p_wishbone_bd_ram_n23125, p_wishbone_bd_ram_n23126,
         p_wishbone_bd_ram_n23127, p_wishbone_bd_ram_n23128,
         p_wishbone_bd_ram_n23129, p_wishbone_bd_ram_n23130,
         p_wishbone_bd_ram_n23131, p_wishbone_bd_ram_n23132,
         p_wishbone_bd_ram_n23133, p_wishbone_bd_ram_n23134,
         p_wishbone_bd_ram_n23135, p_wishbone_bd_ram_n23136,
         p_wishbone_bd_ram_n23137, p_wishbone_bd_ram_n23138,
         p_wishbone_bd_ram_n23139, p_wishbone_bd_ram_n23140,
         p_wishbone_bd_ram_n23141, p_wishbone_bd_ram_n23142,
         p_wishbone_bd_ram_n23143, p_wishbone_bd_ram_n23144,
         p_wishbone_bd_ram_n23145, p_wishbone_bd_ram_n23146,
         p_wishbone_bd_ram_n23147, p_wishbone_bd_ram_n23148,
         p_wishbone_bd_ram_n23149, p_wishbone_bd_ram_n23150,
         p_wishbone_bd_ram_n23151, p_wishbone_bd_ram_n23152,
         p_wishbone_bd_ram_n23153, p_wishbone_bd_ram_n23154,
         p_wishbone_bd_ram_n23155, p_wishbone_bd_ram_n23156,
         p_wishbone_bd_ram_n23157, p_wishbone_bd_ram_n23158,
         p_wishbone_bd_ram_n23159, p_wishbone_bd_ram_n23160,
         p_wishbone_bd_ram_n23161, p_wishbone_bd_ram_n23162,
         p_wishbone_bd_ram_n23163, p_wishbone_bd_ram_n23164,
         p_wishbone_bd_ram_n23165, p_wishbone_bd_ram_n23166,
         p_wishbone_bd_ram_n23167, p_wishbone_bd_ram_n23168,
         p_wishbone_bd_ram_n23169, p_wishbone_bd_ram_n23170,
         p_wishbone_bd_ram_n23171, p_wishbone_bd_ram_n23172,
         p_wishbone_bd_ram_n23173, p_wishbone_bd_ram_n23174,
         p_wishbone_bd_ram_n23175, p_wishbone_bd_ram_n23176,
         p_wishbone_bd_ram_n23177, p_wishbone_bd_ram_n23178,
         p_wishbone_bd_ram_n23179, p_wishbone_bd_ram_n23180,
         p_wishbone_bd_ram_n23181, p_wishbone_bd_ram_n23182,
         p_wishbone_bd_ram_n23183, p_wishbone_bd_ram_n23184,
         p_wishbone_bd_ram_n23185, p_wishbone_bd_ram_n23186,
         p_wishbone_bd_ram_n23187, p_wishbone_bd_ram_n23188,
         p_wishbone_bd_ram_n23189, p_wishbone_bd_ram_n23190,
         p_wishbone_bd_ram_n23191, p_wishbone_bd_ram_n23192,
         p_wishbone_bd_ram_n23193, p_wishbone_bd_ram_n23194,
         p_wishbone_bd_ram_n23195, p_wishbone_bd_ram_n23196,
         p_wishbone_bd_ram_n23197, p_wishbone_bd_ram_n23198,
         p_wishbone_bd_ram_n23199, p_wishbone_bd_ram_n23200,
         p_wishbone_bd_ram_n23201, p_wishbone_bd_ram_n23202,
         p_wishbone_bd_ram_n23203, p_wishbone_bd_ram_n23204,
         p_wishbone_bd_ram_n23205, p_wishbone_bd_ram_n23206,
         p_wishbone_bd_ram_n23207, p_wishbone_bd_ram_n23208,
         p_wishbone_bd_ram_n23209, p_wishbone_bd_ram_n23210,
         p_wishbone_bd_ram_n23211, p_wishbone_bd_ram_n23212,
         p_wishbone_bd_ram_n23213, p_wishbone_bd_ram_n23214,
         p_wishbone_bd_ram_n23215, p_wishbone_bd_ram_n23216,
         p_wishbone_bd_ram_n23217, p_wishbone_bd_ram_n23218,
         p_wishbone_bd_ram_n23219, p_wishbone_bd_ram_n23220,
         p_wishbone_bd_ram_n23221, p_wishbone_bd_ram_n23222,
         p_wishbone_bd_ram_n23223, p_wishbone_bd_ram_n23224,
         p_wishbone_bd_ram_n23225, p_wishbone_bd_ram_n23226,
         p_wishbone_bd_ram_n23227, p_wishbone_bd_ram_n23228,
         p_wishbone_bd_ram_n23229, p_wishbone_bd_ram_n23230,
         p_wishbone_bd_ram_n23231, p_wishbone_bd_ram_n23232,
         p_wishbone_bd_ram_n23233, p_wishbone_bd_ram_n23234,
         p_wishbone_bd_ram_n23235, p_wishbone_bd_ram_n23236,
         p_wishbone_bd_ram_n23237, p_wishbone_bd_ram_n23238,
         p_wishbone_bd_ram_n23239, p_wishbone_bd_ram_n23240,
         p_wishbone_bd_ram_n23241, p_wishbone_bd_ram_n23242,
         p_wishbone_bd_ram_n23243, p_wishbone_bd_ram_n23244,
         p_wishbone_bd_ram_n23245, p_wishbone_bd_ram_n23246,
         p_wishbone_bd_ram_n23247, p_wishbone_bd_ram_n23248,
         p_wishbone_bd_ram_n23249, p_wishbone_bd_ram_n23250,
         p_wishbone_bd_ram_n23251, p_wishbone_bd_ram_n23252,
         p_wishbone_bd_ram_n23253, p_wishbone_bd_ram_n23254,
         p_wishbone_bd_ram_n23255, p_wishbone_bd_ram_n23256,
         p_wishbone_bd_ram_n23257, p_wishbone_bd_ram_n23258,
         p_wishbone_bd_ram_n23259, p_wishbone_bd_ram_n23260,
         p_wishbone_bd_ram_n23261, p_wishbone_bd_ram_n23262,
         p_wishbone_bd_ram_n23263, p_wishbone_bd_ram_n23264,
         p_wishbone_bd_ram_n23265, p_wishbone_bd_ram_n23266,
         p_wishbone_bd_ram_n23267, p_wishbone_bd_ram_n23268,
         p_wishbone_bd_ram_n23269, p_wishbone_bd_ram_n23270,
         p_wishbone_bd_ram_n23271, p_wishbone_bd_ram_n23272,
         p_wishbone_bd_ram_n23273, p_wishbone_bd_ram_n23274,
         p_wishbone_bd_ram_n23275, p_wishbone_bd_ram_n23276,
         p_wishbone_bd_ram_n23277, p_wishbone_bd_ram_n23278,
         p_wishbone_bd_ram_n23279, p_wishbone_bd_ram_n23280,
         p_wishbone_bd_ram_n23281, p_wishbone_bd_ram_n23282,
         p_wishbone_bd_ram_n23283, p_wishbone_bd_ram_n23284,
         p_wishbone_bd_ram_n23285, p_wishbone_bd_ram_n23286,
         p_wishbone_bd_ram_n23287, p_wishbone_bd_ram_n23288,
         p_wishbone_bd_ram_n23289, p_wishbone_bd_ram_n23290,
         p_wishbone_bd_ram_n23291, p_wishbone_bd_ram_n23292,
         p_wishbone_bd_ram_n23293, p_wishbone_bd_ram_n23294,
         p_wishbone_bd_ram_n23295, p_wishbone_bd_ram_n23296,
         p_wishbone_bd_ram_n23297, p_wishbone_bd_ram_n23298,
         p_wishbone_bd_ram_n23299, p_wishbone_bd_ram_n23300,
         p_wishbone_bd_ram_n23301, p_wishbone_bd_ram_n23302,
         p_wishbone_bd_ram_n23303, p_wishbone_bd_ram_n23304,
         p_wishbone_bd_ram_n23305, p_wishbone_bd_ram_n23306,
         p_wishbone_bd_ram_n23307, p_wishbone_bd_ram_n23308,
         p_wishbone_bd_ram_n23309, p_wishbone_bd_ram_n23310,
         p_wishbone_bd_ram_n23311, p_wishbone_bd_ram_n23312,
         p_wishbone_bd_ram_n23313, p_wishbone_bd_ram_n23314,
         p_wishbone_bd_ram_n23315, p_wishbone_bd_ram_n23316,
         p_wishbone_bd_ram_n23317, p_wishbone_bd_ram_n23318,
         p_wishbone_bd_ram_n23319, p_wishbone_bd_ram_n23320,
         p_wishbone_bd_ram_n23321, p_wishbone_bd_ram_n23322,
         p_wishbone_bd_ram_n23323, p_wishbone_bd_ram_n23324,
         p_wishbone_bd_ram_n23325, p_wishbone_bd_ram_n23326,
         p_wishbone_bd_ram_n23327, p_wishbone_bd_ram_n23328,
         p_wishbone_bd_ram_n23329, p_wishbone_bd_ram_n23330,
         p_wishbone_bd_ram_n23331, p_wishbone_bd_ram_n23332,
         p_wishbone_bd_ram_n23333, p_wishbone_bd_ram_n23334,
         p_wishbone_bd_ram_n23335, p_wishbone_bd_ram_n23336,
         p_wishbone_bd_ram_n23337, p_wishbone_bd_ram_n23338,
         p_wishbone_bd_ram_n23339, p_wishbone_bd_ram_n23340,
         p_wishbone_bd_ram_n23341, p_wishbone_bd_ram_n23342,
         p_wishbone_bd_ram_n23343, p_wishbone_bd_ram_n23344,
         p_wishbone_bd_ram_n23345, p_wishbone_bd_ram_n23346,
         p_wishbone_bd_ram_n23347, p_wishbone_bd_ram_n23348,
         p_wishbone_bd_ram_n23349, p_wishbone_bd_ram_n23350,
         p_wishbone_bd_ram_n23351, p_wishbone_bd_ram_n23352,
         p_wishbone_bd_ram_n23353, p_wishbone_bd_ram_n23354,
         p_wishbone_bd_ram_n23355, p_wishbone_bd_ram_n23356,
         p_wishbone_bd_ram_n23357, p_wishbone_bd_ram_n23358,
         p_wishbone_bd_ram_n23359, p_wishbone_bd_ram_n23360,
         p_wishbone_bd_ram_n23361, p_wishbone_bd_ram_n23362,
         p_wishbone_bd_ram_n23363, p_wishbone_bd_ram_n23364,
         p_wishbone_bd_ram_n23365, p_wishbone_bd_ram_n23366,
         p_wishbone_bd_ram_n23367, p_wishbone_bd_ram_n23368,
         p_wishbone_bd_ram_n23369, p_wishbone_bd_ram_n23370,
         p_wishbone_bd_ram_n23371, p_wishbone_bd_ram_n23372,
         p_wishbone_bd_ram_n23373, p_wishbone_bd_ram_n23374,
         p_wishbone_bd_ram_n23375, p_wishbone_bd_ram_n23376,
         p_wishbone_bd_ram_n23377, p_wishbone_bd_ram_n23378,
         p_wishbone_bd_ram_n23379, p_wishbone_bd_ram_n23380,
         p_wishbone_bd_ram_n23381, p_wishbone_bd_ram_n23382,
         p_wishbone_bd_ram_n23383, p_wishbone_bd_ram_n23384,
         p_wishbone_bd_ram_n23385, p_wishbone_bd_ram_n23386,
         p_wishbone_bd_ram_n23387, p_wishbone_bd_ram_n23388,
         p_wishbone_bd_ram_n23389, p_wishbone_bd_ram_n23390,
         p_wishbone_bd_ram_n23391, p_wishbone_bd_ram_n23392,
         p_wishbone_bd_ram_n23393, p_wishbone_bd_ram_n23394,
         p_wishbone_bd_ram_n23395, p_wishbone_bd_ram_n23396,
         p_wishbone_bd_ram_n23397, p_wishbone_bd_ram_n23398,
         p_wishbone_bd_ram_n23399, p_wishbone_bd_ram_n23400,
         p_wishbone_bd_ram_n23401, p_wishbone_bd_ram_n23402,
         p_wishbone_bd_ram_n23403, p_wishbone_bd_ram_n23404,
         p_wishbone_bd_ram_n23405, p_wishbone_bd_ram_n23406,
         p_wishbone_bd_ram_n23407, p_wishbone_bd_ram_n23408,
         p_wishbone_bd_ram_n23409, p_wishbone_bd_ram_n23410,
         p_wishbone_bd_ram_n23411, p_wishbone_bd_ram_n23412,
         p_wishbone_bd_ram_n23413, p_wishbone_bd_ram_n23414,
         p_wishbone_bd_ram_n23415, p_wishbone_bd_ram_n23416,
         p_wishbone_bd_ram_n23417, p_wishbone_bd_ram_n23418,
         p_wishbone_bd_ram_n23419, p_wishbone_bd_ram_n23420,
         p_wishbone_bd_ram_n23421, p_wishbone_bd_ram_n23422,
         p_wishbone_bd_ram_n23423, p_wishbone_bd_ram_n23424,
         p_wishbone_bd_ram_n23425, p_wishbone_bd_ram_n23426,
         p_wishbone_bd_ram_n23427, p_wishbone_bd_ram_n23428,
         p_wishbone_bd_ram_n23429, p_wishbone_bd_ram_n23430,
         p_wishbone_bd_ram_n23431, p_wishbone_bd_ram_n23432,
         p_wishbone_bd_ram_n23433, p_wishbone_bd_ram_n23434,
         p_wishbone_bd_ram_n23435, p_wishbone_bd_ram_n23436,
         p_wishbone_bd_ram_n23437, p_wishbone_bd_ram_n23438,
         p_wishbone_bd_ram_n23439, p_wishbone_bd_ram_n23440,
         p_wishbone_bd_ram_n23441, p_wishbone_bd_ram_n23442,
         p_wishbone_bd_ram_n23443, p_wishbone_bd_ram_n23444,
         p_wishbone_bd_ram_n23445, p_wishbone_bd_ram_n23446,
         p_wishbone_bd_ram_n23447, p_wishbone_bd_ram_n23448,
         p_wishbone_bd_ram_n23449, p_wishbone_bd_ram_n23450,
         p_wishbone_bd_ram_n23451, p_wishbone_bd_ram_n23452,
         p_wishbone_bd_ram_n23453, p_wishbone_bd_ram_n23454,
         p_wishbone_bd_ram_n23455, p_wishbone_bd_ram_n23456,
         p_wishbone_bd_ram_n23457, p_wishbone_bd_ram_n23458,
         p_wishbone_bd_ram_n23459, p_wishbone_bd_ram_n23460,
         p_wishbone_bd_ram_n23461, p_wishbone_bd_ram_n23462,
         p_wishbone_bd_ram_n23463, p_wishbone_bd_ram_n23464,
         p_wishbone_bd_ram_n23465, p_wishbone_bd_ram_n23466,
         p_wishbone_bd_ram_n23467, p_wishbone_bd_ram_n23468,
         p_wishbone_bd_ram_n23469, p_wishbone_bd_ram_n23470,
         p_wishbone_bd_ram_n23471, p_wishbone_bd_ram_n23472,
         p_wishbone_bd_ram_n23473, p_wishbone_bd_ram_n23474,
         p_wishbone_bd_ram_n23475, p_wishbone_bd_ram_n23476,
         p_wishbone_bd_ram_n23477, p_wishbone_bd_ram_n23478,
         p_wishbone_bd_ram_n23479, p_wishbone_bd_ram_n23480,
         p_wishbone_bd_ram_n23481, p_wishbone_bd_ram_n23482,
         p_wishbone_bd_ram_n23483, p_wishbone_bd_ram_n23484,
         p_wishbone_bd_ram_n23485, p_wishbone_bd_ram_n23486,
         p_wishbone_bd_ram_n23487, p_wishbone_bd_ram_n23488,
         p_wishbone_bd_ram_n23489, p_wishbone_bd_ram_n23490,
         p_wishbone_bd_ram_n23491, p_wishbone_bd_ram_n23492,
         p_wishbone_bd_ram_n23493, p_wishbone_bd_ram_n23494,
         p_wishbone_bd_ram_n23495, p_wishbone_bd_ram_n23496,
         p_wishbone_bd_ram_n23497, p_wishbone_bd_ram_n23498,
         p_wishbone_bd_ram_n23499, p_wishbone_bd_ram_n23500,
         p_wishbone_bd_ram_n23501, p_wishbone_bd_ram_n23502,
         p_wishbone_bd_ram_n23503, p_wishbone_bd_ram_n23504,
         p_wishbone_bd_ram_n23505, p_wishbone_bd_ram_n23506,
         p_wishbone_bd_ram_n23507, p_wishbone_bd_ram_n23508,
         p_wishbone_bd_ram_n23509, p_wishbone_bd_ram_n23510,
         p_wishbone_bd_ram_n23511, p_wishbone_bd_ram_n23512,
         p_wishbone_bd_ram_n23513, p_wishbone_bd_ram_n23514,
         p_wishbone_bd_ram_n23515, p_wishbone_bd_ram_n23516,
         p_wishbone_bd_ram_n23517, p_wishbone_bd_ram_n23518,
         p_wishbone_bd_ram_n23519, p_wishbone_bd_ram_n23520,
         p_wishbone_bd_ram_n23521, p_wishbone_bd_ram_n23522,
         p_wishbone_bd_ram_n23523, p_wishbone_bd_ram_n23524,
         p_wishbone_bd_ram_n23525, p_wishbone_bd_ram_n23526,
         p_wishbone_bd_ram_n23527, p_wishbone_bd_ram_n23528,
         p_wishbone_bd_ram_n23529, p_wishbone_bd_ram_n23530,
         p_wishbone_bd_ram_n23531, p_wishbone_bd_ram_n23532,
         p_wishbone_bd_ram_n23533, p_wishbone_bd_ram_n23534,
         p_wishbone_bd_ram_n23535, p_wishbone_bd_ram_n23536,
         p_wishbone_bd_ram_n23537, p_wishbone_bd_ram_n23538,
         p_wishbone_bd_ram_n23539, p_wishbone_bd_ram_n23540,
         p_wishbone_bd_ram_n23541, p_wishbone_bd_ram_n23542,
         p_wishbone_bd_ram_n23543, p_wishbone_bd_ram_n23544,
         p_wishbone_bd_ram_n23545, p_wishbone_bd_ram_n23546,
         p_wishbone_bd_ram_n23547, p_wishbone_bd_ram_n23548,
         p_wishbone_bd_ram_n23549, p_wishbone_bd_ram_n23550,
         p_wishbone_bd_ram_n23551, p_wishbone_bd_ram_n23552,
         p_wishbone_bd_ram_n23553, p_wishbone_bd_ram_n23554,
         p_wishbone_bd_ram_n23555, p_wishbone_bd_ram_n23556,
         p_wishbone_bd_ram_n23557, p_wishbone_bd_ram_n23558,
         p_wishbone_bd_ram_n23559, p_wishbone_bd_ram_n23560,
         p_wishbone_bd_ram_n23561, p_wishbone_bd_ram_n23562,
         p_wishbone_bd_ram_n23563, p_wishbone_bd_ram_n23564,
         p_wishbone_bd_ram_n23565, p_wishbone_bd_ram_n23566,
         p_wishbone_bd_ram_n23567, p_wishbone_bd_ram_n23568,
         p_wishbone_bd_ram_n23569, p_wishbone_bd_ram_n23570,
         p_wishbone_bd_ram_n23571, p_wishbone_bd_ram_n23572,
         p_wishbone_bd_ram_n23573, p_wishbone_bd_ram_n23574,
         p_wishbone_bd_ram_n23575, p_wishbone_bd_ram_n23576,
         p_wishbone_bd_ram_n23577, p_wishbone_bd_ram_n23578,
         p_wishbone_bd_ram_n23579, p_wishbone_bd_ram_n23580,
         p_wishbone_bd_ram_n23581, p_wishbone_bd_ram_n23582,
         p_wishbone_bd_ram_n23583, p_wishbone_bd_ram_n23584,
         p_wishbone_bd_ram_n23585, p_wishbone_bd_ram_n23586,
         p_wishbone_bd_ram_n23587, p_wishbone_bd_ram_n23588,
         p_wishbone_bd_ram_n23589, p_wishbone_bd_ram_n23590,
         p_wishbone_bd_ram_n23591, p_wishbone_bd_ram_n23592,
         p_wishbone_bd_ram_n23593, p_wishbone_bd_ram_n23594,
         p_wishbone_bd_ram_n23595, p_wishbone_bd_ram_n23596,
         p_wishbone_bd_ram_n23597, p_wishbone_bd_ram_n23598,
         p_wishbone_bd_ram_n23599, p_wishbone_bd_ram_n23600,
         p_wishbone_bd_ram_n23601, p_wishbone_bd_ram_n23602,
         p_wishbone_bd_ram_n23603, p_wishbone_bd_ram_n23604,
         p_wishbone_bd_ram_n23605, p_wishbone_bd_ram_n23606,
         p_wishbone_bd_ram_n23607, p_wishbone_bd_ram_n23608,
         p_wishbone_bd_ram_n23609, p_wishbone_bd_ram_n23610,
         p_wishbone_bd_ram_n23611, p_wishbone_bd_ram_n23612,
         p_wishbone_bd_ram_n23613, p_wishbone_bd_ram_n23614,
         p_wishbone_bd_ram_n23615, p_wishbone_bd_ram_n23616,
         p_wishbone_bd_ram_n23617, p_wishbone_bd_ram_n23618,
         p_wishbone_bd_ram_n23619, p_wishbone_bd_ram_n23620,
         p_wishbone_bd_ram_n23621, p_wishbone_bd_ram_n23622,
         p_wishbone_bd_ram_n23623, p_wishbone_bd_ram_n23624,
         p_wishbone_bd_ram_n23625, p_wishbone_bd_ram_n23626,
         p_wishbone_bd_ram_n23627, p_wishbone_bd_ram_n23628,
         p_wishbone_bd_ram_n23629, p_wishbone_bd_ram_n23630,
         p_wishbone_bd_ram_n23631, p_wishbone_bd_ram_n23632,
         p_wishbone_bd_ram_n23633, p_wishbone_bd_ram_n23634,
         p_wishbone_bd_ram_n23635, p_wishbone_bd_ram_n23636,
         p_wishbone_bd_ram_n23637, p_wishbone_bd_ram_n23638,
         p_wishbone_bd_ram_n23639, p_wishbone_bd_ram_n23640,
         p_wishbone_bd_ram_n23641, p_wishbone_bd_ram_n23642,
         p_wishbone_bd_ram_n23643, p_wishbone_bd_ram_n23644,
         p_wishbone_bd_ram_n23645, p_wishbone_bd_ram_n23646,
         p_wishbone_bd_ram_n23647, p_wishbone_bd_ram_n23648,
         p_wishbone_bd_ram_n23649, p_wishbone_bd_ram_n23650,
         p_wishbone_bd_ram_n23651, p_wishbone_bd_ram_n23652,
         p_wishbone_bd_ram_n23653, p_wishbone_bd_ram_n23654,
         p_wishbone_bd_ram_n23655, p_wishbone_bd_ram_n23656,
         p_wishbone_bd_ram_n23657, p_wishbone_bd_ram_n23658,
         p_wishbone_bd_ram_n23659, p_wishbone_bd_ram_n23660,
         p_wishbone_bd_ram_n23661, p_wishbone_bd_ram_n23662,
         p_wishbone_bd_ram_n23663, p_wishbone_bd_ram_n23664,
         p_wishbone_bd_ram_n23665, p_wishbone_bd_ram_n23666,
         p_wishbone_bd_ram_n23667, p_wishbone_bd_ram_n23668,
         p_wishbone_bd_ram_n23669, p_wishbone_bd_ram_n23670,
         p_wishbone_bd_ram_n23671, p_wishbone_bd_ram_n23672,
         p_wishbone_bd_ram_n23673, p_wishbone_bd_ram_n23674,
         p_wishbone_bd_ram_n23675, p_wishbone_bd_ram_n23676,
         p_wishbone_bd_ram_n23677, p_wishbone_bd_ram_n23678,
         p_wishbone_bd_ram_n23679, p_wishbone_bd_ram_n23680,
         p_wishbone_bd_ram_n23681, p_wishbone_bd_ram_n23682,
         p_wishbone_bd_ram_n23683, p_wishbone_bd_ram_n23684,
         p_wishbone_bd_ram_n23685, p_wishbone_bd_ram_n23686,
         p_wishbone_bd_ram_n23687, p_wishbone_bd_ram_n23688,
         p_wishbone_bd_ram_n23689, p_wishbone_bd_ram_n23690,
         p_wishbone_bd_ram_n23691, p_wishbone_bd_ram_n23692,
         p_wishbone_bd_ram_n23693, p_wishbone_bd_ram_n23694,
         p_wishbone_bd_ram_n23695, p_wishbone_bd_ram_n23696,
         p_wishbone_bd_ram_n23697, p_wishbone_bd_ram_n23698,
         p_wishbone_bd_ram_n23699, p_wishbone_bd_ram_n23700,
         p_wishbone_bd_ram_n23701, p_wishbone_bd_ram_n23702,
         p_wishbone_bd_ram_n23703, p_wishbone_bd_ram_n23704,
         p_wishbone_bd_ram_n23705, p_wishbone_bd_ram_n23706,
         p_wishbone_bd_ram_n23707, p_wishbone_bd_ram_n23708,
         p_wishbone_bd_ram_n23709, p_wishbone_bd_ram_n23710,
         p_wishbone_bd_ram_n23711, p_wishbone_bd_ram_n23712,
         p_wishbone_bd_ram_n23713, p_wishbone_bd_ram_n23714,
         p_wishbone_bd_ram_n23715, p_wishbone_bd_ram_n23716,
         p_wishbone_bd_ram_n23717, p_wishbone_bd_ram_n23718,
         p_wishbone_bd_ram_n23719, p_wishbone_bd_ram_n23720,
         p_wishbone_bd_ram_n23721, p_wishbone_bd_ram_n23722,
         p_wishbone_bd_ram_n23723, p_wishbone_bd_ram_n23724,
         p_wishbone_bd_ram_n23725, p_wishbone_bd_ram_n23726,
         p_wishbone_bd_ram_n23727, p_wishbone_bd_ram_n23728,
         p_wishbone_bd_ram_n23729, p_wishbone_bd_ram_n23730,
         p_wishbone_bd_ram_n23731, p_wishbone_bd_ram_n23732,
         p_wishbone_bd_ram_n23733, p_wishbone_bd_ram_n23734,
         p_wishbone_bd_ram_n23735, p_wishbone_bd_ram_n23736,
         p_wishbone_bd_ram_n23737, p_wishbone_bd_ram_n23738,
         p_wishbone_bd_ram_n23739, p_wishbone_bd_ram_n23740,
         p_wishbone_bd_ram_n23741, p_wishbone_bd_ram_n23742,
         p_wishbone_bd_ram_n23743, p_wishbone_bd_ram_n23744,
         p_wishbone_bd_ram_n23745, p_wishbone_bd_ram_n23746,
         p_wishbone_bd_ram_n23747, p_wishbone_bd_ram_n23748,
         p_wishbone_bd_ram_n23749, p_wishbone_bd_ram_n23750,
         p_wishbone_bd_ram_n23751, p_wishbone_bd_ram_n23752,
         p_wishbone_bd_ram_n23753, p_wishbone_bd_ram_n23754,
         p_wishbone_bd_ram_n23755, p_wishbone_bd_ram_n23756,
         p_wishbone_bd_ram_n23757, p_wishbone_bd_ram_n23758,
         p_wishbone_bd_ram_n23759, p_wishbone_bd_ram_n23760,
         p_wishbone_bd_ram_n23761, p_wishbone_bd_ram_n23762,
         p_wishbone_bd_ram_n23763, p_wishbone_bd_ram_n23764,
         p_wishbone_bd_ram_n23765, p_wishbone_bd_ram_n23766,
         p_wishbone_bd_ram_n23767, p_wishbone_bd_ram_n23768,
         p_wishbone_bd_ram_n23769, p_wishbone_bd_ram_n23770,
         p_wishbone_bd_ram_n23771, p_wishbone_bd_ram_n23772,
         p_wishbone_bd_ram_n23773, p_wishbone_bd_ram_n23774,
         p_wishbone_bd_ram_n23775, p_wishbone_bd_ram_n23776,
         p_wishbone_bd_ram_n23777, p_wishbone_bd_ram_n23778,
         p_wishbone_bd_ram_n23779, p_wishbone_bd_ram_n23780,
         p_wishbone_bd_ram_n23781, p_wishbone_bd_ram_n23782,
         p_wishbone_bd_ram_n23783, p_wishbone_bd_ram_n23784,
         p_wishbone_bd_ram_n23785, p_wishbone_bd_ram_n23786,
         p_wishbone_bd_ram_n23787, p_wishbone_bd_ram_n23788,
         p_wishbone_bd_ram_n23789, p_wishbone_bd_ram_n23790,
         p_wishbone_bd_ram_n23791, p_wishbone_bd_ram_n23792,
         p_wishbone_bd_ram_n23793, p_wishbone_bd_ram_n23794,
         p_wishbone_bd_ram_n23795, p_wishbone_bd_ram_n23796,
         p_wishbone_bd_ram_n23797, p_wishbone_bd_ram_n23798,
         p_wishbone_bd_ram_n23799, p_wishbone_bd_ram_n23800,
         p_wishbone_bd_ram_n23801, p_wishbone_bd_ram_n23802,
         p_wishbone_bd_ram_n23803, p_wishbone_bd_ram_n23804,
         p_wishbone_bd_ram_n23805, p_wishbone_bd_ram_n23806,
         p_wishbone_bd_ram_n23807, p_wishbone_bd_ram_n23808,
         p_wishbone_bd_ram_n23809, p_wishbone_bd_ram_n23810,
         p_wishbone_bd_ram_n23811, p_wishbone_bd_ram_n23812,
         p_wishbone_bd_ram_n23813, p_wishbone_bd_ram_n23814,
         p_wishbone_bd_ram_n23815, p_wishbone_bd_ram_n23816,
         p_wishbone_bd_ram_n23817, p_wishbone_bd_ram_n23818,
         p_wishbone_bd_ram_n23819, p_wishbone_bd_ram_n23820,
         p_wishbone_bd_ram_n23821, p_wishbone_bd_ram_n23822,
         p_wishbone_bd_ram_n23823, p_wishbone_bd_ram_n23824,
         p_wishbone_bd_ram_n23825, p_wishbone_bd_ram_n23826,
         p_wishbone_bd_ram_n23827, p_wishbone_bd_ram_n23828,
         p_wishbone_bd_ram_n23829, p_wishbone_bd_ram_n23830,
         p_wishbone_bd_ram_n23831, p_wishbone_bd_ram_n23832,
         p_wishbone_bd_ram_n23833, p_wishbone_bd_ram_n23834,
         p_wishbone_bd_ram_n23835, p_wishbone_bd_ram_n23836,
         p_wishbone_bd_ram_n23837, p_wishbone_bd_ram_n23838,
         p_wishbone_bd_ram_n23839, p_wishbone_bd_ram_n23840,
         p_wishbone_bd_ram_n23841, p_wishbone_bd_ram_n23842,
         p_wishbone_bd_ram_n23843, p_wishbone_bd_ram_n23844,
         p_wishbone_bd_ram_n23845, p_wishbone_bd_ram_n23846,
         p_wishbone_bd_ram_n23847, p_wishbone_bd_ram_n23848,
         p_wishbone_bd_ram_n23849, p_wishbone_bd_ram_n23850,
         p_wishbone_bd_ram_n23851, p_wishbone_bd_ram_n23852,
         p_wishbone_bd_ram_n23853, p_wishbone_bd_ram_n23854,
         p_wishbone_bd_ram_n23855, p_wishbone_bd_ram_n23856,
         p_wishbone_bd_ram_n23857, p_wishbone_bd_ram_n23858,
         p_wishbone_bd_ram_n23859, p_wishbone_bd_ram_n23860,
         p_wishbone_bd_ram_n23861, p_wishbone_bd_ram_n23862,
         p_wishbone_bd_ram_n23863, p_wishbone_bd_ram_n23864,
         p_wishbone_bd_ram_n23865, p_wishbone_bd_ram_n23866,
         p_wishbone_bd_ram_n23867, p_wishbone_bd_ram_n23868,
         p_wishbone_bd_ram_n23869, p_wishbone_bd_ram_n23870,
         p_wishbone_bd_ram_n23871, p_wishbone_bd_ram_n23872,
         p_wishbone_bd_ram_n23873, p_wishbone_bd_ram_n23874,
         p_wishbone_bd_ram_n23875, p_wishbone_bd_ram_n23876,
         p_wishbone_bd_ram_n23877, p_wishbone_bd_ram_n23878,
         p_wishbone_bd_ram_n23879, p_wishbone_bd_ram_n23880,
         p_wishbone_bd_ram_n23881, p_wishbone_bd_ram_n23882,
         p_wishbone_bd_ram_n23883, p_wishbone_bd_ram_n23884,
         p_wishbone_bd_ram_n23885, p_wishbone_bd_ram_n23886,
         p_wishbone_bd_ram_n23887, p_wishbone_bd_ram_n23888,
         p_wishbone_bd_ram_n23889, p_wishbone_bd_ram_n23890,
         p_wishbone_bd_ram_n23891, p_wishbone_bd_ram_n23892,
         p_wishbone_bd_ram_n23893, p_wishbone_bd_ram_n23894,
         p_wishbone_bd_ram_n23895, p_wishbone_bd_ram_n23896,
         p_wishbone_bd_ram_n23897, p_wishbone_bd_ram_n23898,
         p_wishbone_bd_ram_n23899, p_wishbone_bd_ram_n23900,
         p_wishbone_bd_ram_n23901, p_wishbone_bd_ram_n23902,
         p_wishbone_bd_ram_n23903, p_wishbone_bd_ram_n23904,
         p_wishbone_bd_ram_n23905, p_wishbone_bd_ram_n23906,
         p_wishbone_bd_ram_n23907, p_wishbone_bd_ram_n23908,
         p_wishbone_bd_ram_n23909, p_wishbone_bd_ram_n23910,
         p_wishbone_bd_ram_n23911, p_wishbone_bd_ram_n23912,
         p_wishbone_bd_ram_n23913, p_wishbone_bd_ram_n23914,
         p_wishbone_bd_ram_n23915, p_wishbone_bd_ram_n23916,
         p_wishbone_bd_ram_n23917, p_wishbone_bd_ram_n23918,
         p_wishbone_bd_ram_n23919, p_wishbone_bd_ram_n23920,
         p_wishbone_bd_ram_n23921, p_wishbone_bd_ram_n23922,
         p_wishbone_bd_ram_n23923, p_wishbone_bd_ram_n23924,
         p_wishbone_bd_ram_n23925, p_wishbone_bd_ram_n23926,
         p_wishbone_bd_ram_n23927, p_wishbone_bd_ram_n23928,
         p_wishbone_bd_ram_n23929, p_wishbone_bd_ram_n23930,
         p_wishbone_bd_ram_n23931, p_wishbone_bd_ram_n23932,
         p_wishbone_bd_ram_n23933, p_wishbone_bd_ram_n23934,
         p_wishbone_bd_ram_n23935, p_wishbone_bd_ram_n23936,
         p_wishbone_bd_ram_n23937, p_wishbone_bd_ram_n23938,
         p_wishbone_bd_ram_n23939, p_wishbone_bd_ram_n23940,
         p_wishbone_bd_ram_n23941, p_wishbone_bd_ram_n23942,
         p_wishbone_bd_ram_n23943, p_wishbone_bd_ram_n23944,
         p_wishbone_bd_ram_n23945, p_wishbone_bd_ram_n23946,
         p_wishbone_bd_ram_n23947, p_wishbone_bd_ram_n23948,
         p_wishbone_bd_ram_n23949, p_wishbone_bd_ram_n23950,
         p_wishbone_bd_ram_n23951, p_wishbone_bd_ram_n23952,
         p_wishbone_bd_ram_n23953, p_wishbone_bd_ram_n23954,
         p_wishbone_bd_ram_n23955, p_wishbone_bd_ram_n23956,
         p_wishbone_bd_ram_n23957, p_wishbone_bd_ram_n23958,
         p_wishbone_bd_ram_n23959, p_wishbone_bd_ram_n23960,
         p_wishbone_bd_ram_n23961, p_wishbone_bd_ram_n23962,
         p_wishbone_bd_ram_n23963, p_wishbone_bd_ram_n23964,
         p_wishbone_bd_ram_n23965, p_wishbone_bd_ram_n23966,
         p_wishbone_bd_ram_n23967, p_wishbone_bd_ram_n23968,
         p_wishbone_bd_ram_n23969, p_wishbone_bd_ram_n23970,
         p_wishbone_bd_ram_n23971, p_wishbone_bd_ram_n23972,
         p_wishbone_bd_ram_n23973, p_wishbone_bd_ram_n23974,
         p_wishbone_bd_ram_n23975, p_wishbone_bd_ram_n23976,
         p_wishbone_bd_ram_n23977, p_wishbone_bd_ram_n23978,
         p_wishbone_bd_ram_n23979, p_wishbone_bd_ram_n23980,
         p_wishbone_bd_ram_n23981, p_wishbone_bd_ram_n23982,
         p_wishbone_bd_ram_n23983, p_wishbone_bd_ram_n23984,
         p_wishbone_bd_ram_n23985, p_wishbone_bd_ram_n23986,
         p_wishbone_bd_ram_n23987, p_wishbone_bd_ram_n23988,
         p_wishbone_bd_ram_n23989, p_wishbone_bd_ram_n23990,
         p_wishbone_bd_ram_n23991, p_wishbone_bd_ram_n23992,
         p_wishbone_bd_ram_n23993, p_wishbone_bd_ram_n23994,
         p_wishbone_bd_ram_n23995, p_wishbone_bd_ram_n23996,
         p_wishbone_bd_ram_n23997, p_wishbone_bd_ram_n23998,
         p_wishbone_bd_ram_n23999, p_wishbone_bd_ram_n24000,
         p_wishbone_bd_ram_n24001, p_wishbone_bd_ram_n24002,
         p_wishbone_bd_ram_n24003, p_wishbone_bd_ram_n24004,
         p_wishbone_bd_ram_n24005, p_wishbone_bd_ram_n24006,
         p_wishbone_bd_ram_n24007, p_wishbone_bd_ram_n24008,
         p_wishbone_bd_ram_n24009, p_wishbone_bd_ram_n24010,
         p_wishbone_bd_ram_n24011, p_wishbone_bd_ram_n24012,
         p_wishbone_bd_ram_n24013, p_wishbone_bd_ram_n24014,
         p_wishbone_bd_ram_n24015, p_wishbone_bd_ram_n24016,
         p_wishbone_bd_ram_n24017, p_wishbone_bd_ram_n24018,
         p_wishbone_bd_ram_n24019, p_wishbone_bd_ram_n24020,
         p_wishbone_bd_ram_n24021, p_wishbone_bd_ram_n24022,
         p_wishbone_bd_ram_n24023, p_wishbone_bd_ram_n24024,
         p_wishbone_bd_ram_n24025, p_wishbone_bd_ram_n24026,
         p_wishbone_bd_ram_n24027, p_wishbone_bd_ram_n24028,
         p_wishbone_bd_ram_n24029, p_wishbone_bd_ram_n24030,
         p_wishbone_bd_ram_n24031, p_wishbone_bd_ram_n24032,
         p_wishbone_bd_ram_n24033, p_wishbone_bd_ram_n24034,
         p_wishbone_bd_ram_n24035, p_wishbone_bd_ram_n24036,
         p_wishbone_bd_ram_n24037, p_wishbone_bd_ram_n24038,
         p_wishbone_bd_ram_n24039, p_wishbone_bd_ram_n24040,
         p_wishbone_bd_ram_n24041, p_wishbone_bd_ram_n24042,
         p_wishbone_bd_ram_n24043, p_wishbone_bd_ram_n24044,
         p_wishbone_bd_ram_n24045, p_wishbone_bd_ram_n24046,
         p_wishbone_bd_ram_n24047, p_wishbone_bd_ram_n24048,
         p_wishbone_bd_ram_n24049, p_wishbone_bd_ram_n24050,
         p_wishbone_bd_ram_n24051, p_wishbone_bd_ram_n24052,
         p_wishbone_bd_ram_n24053, p_wishbone_bd_ram_n24054,
         p_wishbone_bd_ram_n24055, p_wishbone_bd_ram_n24056,
         p_wishbone_bd_ram_n24057, p_wishbone_bd_ram_n24058,
         p_wishbone_bd_ram_n24059, p_wishbone_bd_ram_n24060,
         p_wishbone_bd_ram_n24061, p_wishbone_bd_ram_n24062,
         p_wishbone_bd_ram_n24063, p_wishbone_bd_ram_n24064,
         p_wishbone_bd_ram_n24065, p_wishbone_bd_ram_n24066,
         p_wishbone_bd_ram_n24067, p_wishbone_bd_ram_n24068,
         p_wishbone_bd_ram_n24069, p_wishbone_bd_ram_n24070,
         p_wishbone_bd_ram_n24071, p_wishbone_bd_ram_n24072,
         p_wishbone_bd_ram_n24073, p_wishbone_bd_ram_n24074,
         p_wishbone_bd_ram_n24075, p_wishbone_bd_ram_n24076,
         p_wishbone_bd_ram_n24077, p_wishbone_bd_ram_n24078,
         p_wishbone_bd_ram_n24079, p_wishbone_bd_ram_n24080,
         p_wishbone_bd_ram_n24081, p_wishbone_bd_ram_n24082,
         p_wishbone_bd_ram_n24083, p_wishbone_bd_ram_n24084,
         p_wishbone_bd_ram_n24085, p_wishbone_bd_ram_n24086,
         p_wishbone_bd_ram_n24087, p_wishbone_bd_ram_n24088,
         p_wishbone_bd_ram_n24089, p_wishbone_bd_ram_n24090,
         p_wishbone_bd_ram_n24091, p_wishbone_bd_ram_n24092,
         p_wishbone_bd_ram_n24093, p_wishbone_bd_ram_n24094,
         p_wishbone_bd_ram_n24095, p_wishbone_bd_ram_n24096,
         p_wishbone_bd_ram_n24097, p_wishbone_bd_ram_n24098,
         p_wishbone_bd_ram_n24099, p_wishbone_bd_ram_n24100,
         p_wishbone_bd_ram_n24101, p_wishbone_bd_ram_n24102,
         p_wishbone_bd_ram_n24103, p_wishbone_bd_ram_n24104,
         p_wishbone_bd_ram_n24105, p_wishbone_bd_ram_n24106,
         p_wishbone_bd_ram_n24107, p_wishbone_bd_ram_n24108,
         p_wishbone_bd_ram_n24109, p_wishbone_bd_ram_n24110,
         p_wishbone_bd_ram_n24111, p_wishbone_bd_ram_n24112,
         p_wishbone_bd_ram_n24113, p_wishbone_bd_ram_n24114,
         p_wishbone_bd_ram_n24115, p_wishbone_bd_ram_n24116,
         p_wishbone_bd_ram_n24117, p_wishbone_bd_ram_n24118,
         p_wishbone_bd_ram_n24119, p_wishbone_bd_ram_n24120,
         p_wishbone_bd_ram_n24121, p_wishbone_bd_ram_n24122,
         p_wishbone_bd_ram_n24123, p_wishbone_bd_ram_n24124,
         p_wishbone_bd_ram_n24125, p_wishbone_bd_ram_n24126,
         p_wishbone_bd_ram_n24127, p_wishbone_bd_ram_n24128,
         p_wishbone_bd_ram_n24129, p_wishbone_bd_ram_n24130,
         p_wishbone_bd_ram_n24131, p_wishbone_bd_ram_n24132,
         p_wishbone_bd_ram_n24133, p_wishbone_bd_ram_n24134,
         p_wishbone_bd_ram_n24135, p_wishbone_bd_ram_n24136,
         p_wishbone_bd_ram_n24137, p_wishbone_bd_ram_n24138,
         p_wishbone_bd_ram_n24139, p_wishbone_bd_ram_n24140,
         p_wishbone_bd_ram_n24141, p_wishbone_bd_ram_n24142,
         p_wishbone_bd_ram_n24143, p_wishbone_bd_ram_n24144,
         p_wishbone_bd_ram_n24145, p_wishbone_bd_ram_n24146,
         p_wishbone_bd_ram_n24147, p_wishbone_bd_ram_n24148,
         p_wishbone_bd_ram_n24149, p_wishbone_bd_ram_n24150,
         p_wishbone_bd_ram_n24151, p_wishbone_bd_ram_n24152,
         p_wishbone_bd_ram_n24153, p_wishbone_bd_ram_n24154,
         p_wishbone_bd_ram_n24155, p_wishbone_bd_ram_n24156,
         p_wishbone_bd_ram_n24157, p_wishbone_bd_ram_n24158,
         p_wishbone_bd_ram_n24159, p_wishbone_bd_ram_n24160,
         p_wishbone_bd_ram_n24161, p_wishbone_bd_ram_n24162,
         p_wishbone_bd_ram_n24163, p_wishbone_bd_ram_n24164,
         p_wishbone_bd_ram_n24165, p_wishbone_bd_ram_n24166,
         p_wishbone_bd_ram_n24167, p_wishbone_bd_ram_n24168,
         p_wishbone_bd_ram_n24169, p_wishbone_bd_ram_n24170,
         p_wishbone_bd_ram_n24171, p_wishbone_bd_ram_n24172,
         p_wishbone_bd_ram_n24173, p_wishbone_bd_ram_n24174,
         p_wishbone_bd_ram_n24175, p_wishbone_bd_ram_n24176,
         p_wishbone_bd_ram_n24177, p_wishbone_bd_ram_n24178,
         p_wishbone_bd_ram_n24179, p_wishbone_bd_ram_n24180,
         p_wishbone_bd_ram_n24181, p_wishbone_bd_ram_n24182,
         p_wishbone_bd_ram_n24183, p_wishbone_bd_ram_n24184,
         p_wishbone_bd_ram_n24185, p_wishbone_bd_ram_n24186,
         p_wishbone_bd_ram_n24187, p_wishbone_bd_ram_n24188,
         p_wishbone_bd_ram_n24189, p_wishbone_bd_ram_n24190,
         p_wishbone_bd_ram_n24191, p_wishbone_bd_ram_n24192,
         p_wishbone_bd_ram_n24193, p_wishbone_bd_ram_n24194,
         p_wishbone_bd_ram_n24195, p_wishbone_bd_ram_n24196,
         p_wishbone_bd_ram_n24197, p_wishbone_bd_ram_n24198,
         p_wishbone_bd_ram_n24199, p_wishbone_bd_ram_n24200,
         p_wishbone_bd_ram_n24201, p_wishbone_bd_ram_n24202,
         p_wishbone_bd_ram_n24203, p_wishbone_bd_ram_n24204,
         p_wishbone_bd_ram_n24205, p_wishbone_bd_ram_n24206,
         p_wishbone_bd_ram_n24207, p_wishbone_bd_ram_n24208,
         p_wishbone_bd_ram_n24209, p_wishbone_bd_ram_n24210,
         p_wishbone_bd_ram_n24211, p_wishbone_bd_ram_n24212,
         p_wishbone_bd_ram_n24213, p_wishbone_bd_ram_n24214,
         p_wishbone_bd_ram_n24215, p_wishbone_bd_ram_n24216,
         p_wishbone_bd_ram_n24217, p_wishbone_bd_ram_n24218,
         p_wishbone_bd_ram_n24219, p_wishbone_bd_ram_n24220,
         p_wishbone_bd_ram_n24221, p_wishbone_bd_ram_n24222,
         p_wishbone_bd_ram_n24223, p_wishbone_bd_ram_n24224,
         p_wishbone_bd_ram_n24225, p_wishbone_bd_ram_n24226,
         p_wishbone_bd_ram_n24227, p_wishbone_bd_ram_n24228,
         p_wishbone_bd_ram_n24229, p_wishbone_bd_ram_n24230,
         p_wishbone_bd_ram_n24231, p_wishbone_bd_ram_n24232,
         p_wishbone_bd_ram_n24233, p_wishbone_bd_ram_n24234,
         p_wishbone_bd_ram_n24235, p_wishbone_bd_ram_n24236,
         p_wishbone_bd_ram_n24237, p_wishbone_bd_ram_n24238,
         p_wishbone_bd_ram_n24239, p_wishbone_bd_ram_n24240,
         p_wishbone_bd_ram_n24241, p_wishbone_bd_ram_n24242,
         p_wishbone_bd_ram_n24243, p_wishbone_bd_ram_n24244,
         p_wishbone_bd_ram_n24245, p_wishbone_bd_ram_n24246,
         p_wishbone_bd_ram_n24247, p_wishbone_bd_ram_n24248,
         p_wishbone_bd_ram_n24249, p_wishbone_bd_ram_n24250,
         p_wishbone_bd_ram_n24251, p_wishbone_bd_ram_n24252,
         p_wishbone_bd_ram_n24253, p_wishbone_bd_ram_n24254,
         p_wishbone_bd_ram_n24255, p_wishbone_bd_ram_n24256,
         p_wishbone_bd_ram_n24257, p_wishbone_bd_ram_n24258,
         p_wishbone_bd_ram_n24259, p_wishbone_bd_ram_n24260,
         p_wishbone_bd_ram_n24261, p_wishbone_bd_ram_n24262,
         p_wishbone_bd_ram_n24263, p_wishbone_bd_ram_n24264,
         p_wishbone_bd_ram_n24265, p_wishbone_bd_ram_n24266,
         p_wishbone_bd_ram_n24267, p_wishbone_bd_ram_n24268,
         p_wishbone_bd_ram_n24269, p_wishbone_bd_ram_n24270,
         p_wishbone_bd_ram_n24271, p_wishbone_bd_ram_n24272,
         p_wishbone_bd_ram_n24273, p_wishbone_bd_ram_n24274,
         p_wishbone_bd_ram_n24275, p_wishbone_bd_ram_n24276,
         p_wishbone_bd_ram_n24277, p_wishbone_bd_ram_n24278,
         p_wishbone_bd_ram_n24279, p_wishbone_bd_ram_n24280,
         p_wishbone_bd_ram_n24281, p_wishbone_bd_ram_n24282,
         p_wishbone_bd_ram_n24283, p_wishbone_bd_ram_n24284,
         p_wishbone_bd_ram_n24285, p_wishbone_bd_ram_n24286,
         p_wishbone_bd_ram_n24287, p_wishbone_bd_ram_n24288,
         p_wishbone_bd_ram_n24289, p_wishbone_bd_ram_n24290,
         p_wishbone_bd_ram_n24291, p_wishbone_bd_ram_n24292,
         p_wishbone_bd_ram_n24293, p_wishbone_bd_ram_n24294,
         p_wishbone_bd_ram_n24295, p_wishbone_bd_ram_n24296,
         p_wishbone_bd_ram_n24297, p_wishbone_bd_ram_n24298,
         p_wishbone_bd_ram_n24299, p_wishbone_bd_ram_n24300,
         p_wishbone_bd_ram_n24301, p_wishbone_bd_ram_n24302,
         p_wishbone_bd_ram_n24303, p_wishbone_bd_ram_n24304,
         p_wishbone_bd_ram_n24305, p_wishbone_bd_ram_n24306,
         p_wishbone_bd_ram_n24307, p_wishbone_bd_ram_n24308,
         p_wishbone_bd_ram_n24309, p_wishbone_bd_ram_n24310,
         p_wishbone_bd_ram_n24311, p_wishbone_bd_ram_n24312,
         p_wishbone_bd_ram_n24313, p_wishbone_bd_ram_n24314,
         p_wishbone_bd_ram_n24315, p_wishbone_bd_ram_n24316,
         p_wishbone_bd_ram_n24317, p_wishbone_bd_ram_n24318,
         p_wishbone_bd_ram_n24319, p_wishbone_bd_ram_n24320,
         p_wishbone_bd_ram_n24321, p_wishbone_bd_ram_n24322,
         p_wishbone_bd_ram_n24323, p_wishbone_bd_ram_n24324,
         p_wishbone_bd_ram_n24325, p_wishbone_bd_ram_n24326,
         p_wishbone_bd_ram_n24327, p_wishbone_bd_ram_n24328,
         p_wishbone_bd_ram_n24329, p_wishbone_bd_ram_n24330,
         p_wishbone_bd_ram_n24331, p_wishbone_bd_ram_n24332,
         p_wishbone_bd_ram_n24333, p_wishbone_bd_ram_n24334,
         p_wishbone_bd_ram_n24335, p_wishbone_bd_ram_n24336,
         p_wishbone_bd_ram_n24337, p_wishbone_bd_ram_n24338,
         p_wishbone_bd_ram_n24339, p_wishbone_bd_ram_n24340,
         p_wishbone_bd_ram_n24341, p_wishbone_bd_ram_n24342,
         p_wishbone_bd_ram_n24343, p_wishbone_bd_ram_n24344,
         p_wishbone_bd_ram_n24345, p_wishbone_bd_ram_n24346,
         p_wishbone_bd_ram_n24347, p_wishbone_bd_ram_n24348,
         p_wishbone_bd_ram_n24349, p_wishbone_bd_ram_n24350,
         p_wishbone_bd_ram_n24351, p_wishbone_bd_ram_n24352,
         p_wishbone_bd_ram_n24353, p_wishbone_bd_ram_n24354,
         p_wishbone_bd_ram_n24355, p_wishbone_bd_ram_n24356,
         p_wishbone_bd_ram_n24357, p_wishbone_bd_ram_n24358,
         p_wishbone_bd_ram_n24359, p_wishbone_bd_ram_n24360,
         p_wishbone_bd_ram_n24361, p_wishbone_bd_ram_n24362,
         p_wishbone_bd_ram_n24363, p_wishbone_bd_ram_n24364,
         p_wishbone_bd_ram_n24365, p_wishbone_bd_ram_n24366,
         p_wishbone_bd_ram_n24367, p_wishbone_bd_ram_n24368,
         p_wishbone_bd_ram_n24369, p_wishbone_bd_ram_n24370,
         p_wishbone_bd_ram_n24371, p_wishbone_bd_ram_n24372,
         p_wishbone_bd_ram_n24373, p_wishbone_bd_ram_n24374,
         p_wishbone_bd_ram_n24375, p_wishbone_bd_ram_n24376,
         p_wishbone_bd_ram_n24377, p_wishbone_bd_ram_n24378,
         p_wishbone_bd_ram_n24379, p_wishbone_bd_ram_n24380,
         p_wishbone_bd_ram_n24381, p_wishbone_bd_ram_n24382,
         p_wishbone_bd_ram_n24383, p_wishbone_bd_ram_n24384,
         p_wishbone_bd_ram_n24385, p_wishbone_bd_ram_n24386,
         p_wishbone_bd_ram_n24387, p_wishbone_bd_ram_n24388,
         p_wishbone_bd_ram_n24389, p_wishbone_bd_ram_n24390,
         p_wishbone_bd_ram_n24391, p_wishbone_bd_ram_n24392,
         p_wishbone_bd_ram_n24393, p_wishbone_bd_ram_n24394,
         p_wishbone_bd_ram_n24395, p_wishbone_bd_ram_n24396,
         p_wishbone_bd_ram_n24397, p_wishbone_bd_ram_n24398,
         p_wishbone_bd_ram_n24399, p_wishbone_bd_ram_n24400,
         p_wishbone_bd_ram_n24401, p_wishbone_bd_ram_n24402,
         p_wishbone_bd_ram_n24403, p_wishbone_bd_ram_n24404,
         p_wishbone_bd_ram_n24405, p_wishbone_bd_ram_n24406,
         p_wishbone_bd_ram_n24407, p_wishbone_bd_ram_n24408,
         p_wishbone_bd_ram_n24409, p_wishbone_bd_ram_n24410,
         p_wishbone_bd_ram_n24411, p_wishbone_bd_ram_n24412,
         p_wishbone_bd_ram_n24413, p_wishbone_bd_ram_n24414,
         p_wishbone_bd_ram_n24415, p_wishbone_bd_ram_n24416,
         p_wishbone_bd_ram_n24417, p_wishbone_bd_ram_n24418,
         p_wishbone_bd_ram_n24419, p_wishbone_bd_ram_n24420,
         p_wishbone_bd_ram_n24421, p_wishbone_bd_ram_n24422,
         p_wishbone_bd_ram_n24423, p_wishbone_bd_ram_n24424,
         p_wishbone_bd_ram_n24425, p_wishbone_bd_ram_n24426,
         p_wishbone_bd_ram_n24427, p_wishbone_bd_ram_n24428,
         p_wishbone_bd_ram_n24429, p_wishbone_bd_ram_n24430,
         p_wishbone_bd_ram_n24431, p_wishbone_bd_ram_n24432,
         p_wishbone_bd_ram_n24433, p_wishbone_bd_ram_n24434,
         p_wishbone_bd_ram_n24435, p_wishbone_bd_ram_n24436,
         p_wishbone_bd_ram_n24437, p_wishbone_bd_ram_n24438,
         p_wishbone_bd_ram_n24439, p_wishbone_bd_ram_n24440,
         p_wishbone_bd_ram_n24441, p_wishbone_bd_ram_n24442,
         p_wishbone_bd_ram_n24443, p_wishbone_bd_ram_n24444,
         p_wishbone_bd_ram_n24445, p_wishbone_bd_ram_n24446,
         p_wishbone_bd_ram_n24447, p_wishbone_bd_ram_n24448,
         p_wishbone_bd_ram_n24449, p_wishbone_bd_ram_n24450,
         p_wishbone_bd_ram_n24451, p_wishbone_bd_ram_n24452,
         p_wishbone_bd_ram_n24453, p_wishbone_bd_ram_n24454,
         p_wishbone_bd_ram_n24455, p_wishbone_bd_ram_n24456,
         p_wishbone_bd_ram_n24457, p_wishbone_bd_ram_n24458,
         p_wishbone_bd_ram_n24459, p_wishbone_bd_ram_n24460,
         p_wishbone_bd_ram_n24461, p_wishbone_bd_ram_n24462,
         p_wishbone_bd_ram_n24463, p_wishbone_bd_ram_n24464,
         p_wishbone_bd_ram_n24465, p_wishbone_bd_ram_n24466,
         p_wishbone_bd_ram_n24467, p_wishbone_bd_ram_n24468,
         p_wishbone_bd_ram_n24469, p_wishbone_bd_ram_n24470,
         p_wishbone_bd_ram_n24471, p_wishbone_bd_ram_n24472,
         p_wishbone_bd_ram_n24473, p_wishbone_bd_ram_n24474,
         p_wishbone_bd_ram_n24475, p_wishbone_bd_ram_n24476,
         p_wishbone_bd_ram_n24477, p_wishbone_bd_ram_n24478,
         p_wishbone_bd_ram_n24479, p_wishbone_bd_ram_n24480,
         p_wishbone_bd_ram_n24481, p_wishbone_bd_ram_n24482,
         p_wishbone_bd_ram_n24483, p_wishbone_bd_ram_n24484,
         p_wishbone_bd_ram_n24485, p_wishbone_bd_ram_n24486,
         p_wishbone_bd_ram_n24487, p_wishbone_bd_ram_n24488,
         p_wishbone_bd_ram_n24489, p_wishbone_bd_ram_n24490,
         p_wishbone_bd_ram_n24491, p_wishbone_bd_ram_n24492,
         p_wishbone_bd_ram_n24493, p_wishbone_bd_ram_n24494,
         p_wishbone_bd_ram_n24495, p_wishbone_bd_ram_n24496,
         p_wishbone_bd_ram_n24497, p_wishbone_bd_ram_n24498,
         p_wishbone_bd_ram_n24499, p_wishbone_bd_ram_n24500,
         p_wishbone_bd_ram_n24501, p_wishbone_bd_ram_n24502,
         p_wishbone_bd_ram_n24503, p_wishbone_bd_ram_n24504,
         p_wishbone_bd_ram_n24505, p_wishbone_bd_ram_n24506,
         p_wishbone_bd_ram_n24507, p_wishbone_bd_ram_n24508,
         p_wishbone_bd_ram_n24509, p_wishbone_bd_ram_n24510,
         p_wishbone_bd_ram_n24511, p_wishbone_bd_ram_n24512,
         p_wishbone_bd_ram_n24513, p_wishbone_bd_ram_n24514,
         p_wishbone_bd_ram_n24515, p_wishbone_bd_ram_n24516,
         p_wishbone_bd_ram_n24517, p_wishbone_bd_ram_n24518,
         p_wishbone_bd_ram_n24519, p_wishbone_bd_ram_n24520,
         p_wishbone_bd_ram_n24521, p_wishbone_bd_ram_n24522,
         p_wishbone_bd_ram_n24523, p_wishbone_bd_ram_n24524,
         p_wishbone_bd_ram_n24525, p_wishbone_bd_ram_n24526,
         p_wishbone_bd_ram_n24527, p_wishbone_bd_ram_n24528,
         p_wishbone_bd_ram_n24529, p_wishbone_bd_ram_n24530,
         p_wishbone_bd_ram_n24531, p_wishbone_bd_ram_n24532,
         p_wishbone_bd_ram_n24533, p_wishbone_bd_ram_n24534,
         p_wishbone_bd_ram_n24535, p_wishbone_bd_ram_n24536,
         p_wishbone_bd_ram_n24537, p_wishbone_bd_ram_n24538,
         p_wishbone_bd_ram_n24539, p_wishbone_bd_ram_n24540,
         p_wishbone_bd_ram_n24541, p_wishbone_bd_ram_n24542,
         p_wishbone_bd_ram_n24543, p_wishbone_bd_ram_n24544,
         p_wishbone_bd_ram_n24545, p_wishbone_bd_ram_n24546,
         p_wishbone_bd_ram_n24547, p_wishbone_bd_ram_n24548,
         p_wishbone_bd_ram_n24549, p_wishbone_bd_ram_n24550,
         p_wishbone_bd_ram_n24551, p_wishbone_bd_ram_n24552,
         p_wishbone_bd_ram_n24553, p_wishbone_bd_ram_n24554,
         p_wishbone_bd_ram_n24555, p_wishbone_bd_ram_n24556,
         p_wishbone_bd_ram_n24557, p_wishbone_bd_ram_n24558,
         p_wishbone_bd_ram_n24559, p_wishbone_bd_ram_n24560,
         p_wishbone_bd_ram_n24561, p_wishbone_bd_ram_n24562,
         p_wishbone_bd_ram_n24563, p_wishbone_bd_ram_n24564,
         p_wishbone_bd_ram_n24565, p_wishbone_bd_ram_n24566,
         p_wishbone_bd_ram_n24567, p_wishbone_bd_ram_n24568,
         p_wishbone_bd_ram_n24569, p_wishbone_bd_ram_n24570,
         p_wishbone_bd_ram_n24571, p_wishbone_bd_ram_n24572,
         p_wishbone_bd_ram_n24573, p_wishbone_bd_ram_n24574,
         p_wishbone_bd_ram_n24575, p_wishbone_bd_ram_n24576,
         p_wishbone_bd_ram_n24577, p_wishbone_bd_ram_n24578,
         p_wishbone_bd_ram_n24579, p_wishbone_bd_ram_n24580,
         p_wishbone_bd_ram_n24581, p_wishbone_bd_ram_n24582,
         p_wishbone_bd_ram_n24583, p_wishbone_bd_ram_n24584,
         p_wishbone_bd_ram_n24585, p_wishbone_bd_ram_n24586,
         p_wishbone_bd_ram_n24587, p_wishbone_bd_ram_n24588,
         p_wishbone_bd_ram_n24589, p_wishbone_bd_ram_n24590,
         p_wishbone_bd_ram_n24591, p_wishbone_bd_ram_n24592,
         p_wishbone_bd_ram_n24593, p_wishbone_bd_ram_n24594,
         p_wishbone_bd_ram_n24595, p_wishbone_bd_ram_n24596,
         p_wishbone_bd_ram_n24597, p_wishbone_bd_ram_n24598,
         p_wishbone_bd_ram_n24599, p_wishbone_bd_ram_n24600,
         p_wishbone_bd_ram_n24601, p_wishbone_bd_ram_n24602,
         p_wishbone_bd_ram_n24603, p_wishbone_bd_ram_n24604,
         p_wishbone_bd_ram_n24605, p_wishbone_bd_ram_n24606,
         p_wishbone_bd_ram_n24607, p_wishbone_bd_ram_n24608,
         p_wishbone_bd_ram_n24609, p_wishbone_bd_ram_n24610,
         p_wishbone_bd_ram_n24611, p_wishbone_bd_ram_n24612,
         p_wishbone_bd_ram_n24613, p_wishbone_bd_ram_n24614,
         p_wishbone_bd_ram_n24615, p_wishbone_bd_ram_n24616,
         p_wishbone_bd_ram_n24617, p_wishbone_bd_ram_n24618,
         p_wishbone_bd_ram_n24619, p_wishbone_bd_ram_n24620,
         p_wishbone_bd_ram_n24621, p_wishbone_bd_ram_n24622,
         p_wishbone_bd_ram_n24623, p_wishbone_bd_ram_n24624,
         p_wishbone_bd_ram_n24625, p_wishbone_bd_ram_n24626,
         p_wishbone_bd_ram_n24627, p_wishbone_bd_ram_n24628,
         p_wishbone_bd_ram_n24629, p_wishbone_bd_ram_n24630,
         p_wishbone_bd_ram_n24631, p_wishbone_bd_ram_n24632,
         p_wishbone_bd_ram_n24633, p_wishbone_bd_ram_n24634,
         p_wishbone_bd_ram_n24635, p_wishbone_bd_ram_n24636,
         p_wishbone_bd_ram_n24637, p_wishbone_bd_ram_n24638,
         p_wishbone_bd_ram_n24639, p_wishbone_bd_ram_n24640,
         p_wishbone_bd_ram_n24641, p_wishbone_bd_ram_n24642,
         p_wishbone_bd_ram_n24643, p_wishbone_bd_ram_n24644,
         p_wishbone_bd_ram_n24645, p_wishbone_bd_ram_n24646,
         p_wishbone_bd_ram_n24647, p_wishbone_bd_ram_n24648,
         p_wishbone_bd_ram_n24649, p_wishbone_bd_ram_n24650,
         p_wishbone_bd_ram_n24651, p_wishbone_bd_ram_n24652,
         p_wishbone_bd_ram_n24653, p_wishbone_bd_ram_n24654,
         p_wishbone_bd_ram_n24655, p_wishbone_bd_ram_n24656,
         p_wishbone_bd_ram_n24657, p_wishbone_bd_ram_n24658,
         p_wishbone_bd_ram_n24659, p_wishbone_bd_ram_n24660,
         p_wishbone_bd_ram_n24661, p_wishbone_bd_ram_n24662,
         p_wishbone_bd_ram_n24663, p_wishbone_bd_ram_n24664,
         p_wishbone_bd_ram_n24665, p_wishbone_bd_ram_n24666,
         p_wishbone_bd_ram_n24667, p_wishbone_bd_ram_n24668,
         p_wishbone_bd_ram_n24669, p_wishbone_bd_ram_n24670,
         p_wishbone_bd_ram_n24671, p_wishbone_bd_ram_n24672,
         p_wishbone_bd_ram_n24673, p_wishbone_bd_ram_n24674,
         p_wishbone_bd_ram_n24675, p_wishbone_bd_ram_n24676,
         p_wishbone_bd_ram_n24677, p_wishbone_bd_ram_n24678,
         p_wishbone_bd_ram_n24679, p_wishbone_bd_ram_n24680,
         p_wishbone_bd_ram_n24681, p_wishbone_bd_ram_n24682,
         p_wishbone_bd_ram_n24683, p_wishbone_bd_ram_n24684,
         p_wishbone_bd_ram_n24685, p_wishbone_bd_ram_n24686,
         p_wishbone_bd_ram_n24687, p_wishbone_bd_ram_n24688,
         p_wishbone_bd_ram_n24689, p_wishbone_bd_ram_n24690,
         p_wishbone_bd_ram_n24691, p_wishbone_bd_ram_n24692,
         p_wishbone_bd_ram_n24693, p_wishbone_bd_ram_n24694,
         p_wishbone_bd_ram_n24695, p_wishbone_bd_ram_n24696,
         p_wishbone_bd_ram_n24697, p_wishbone_bd_ram_n24698,
         p_wishbone_bd_ram_n24699, p_wishbone_bd_ram_n24700,
         p_wishbone_bd_ram_n24701, p_wishbone_bd_ram_n24702,
         p_wishbone_bd_ram_n24703, p_wishbone_bd_ram_n24704,
         p_wishbone_bd_ram_n24705, p_wishbone_bd_ram_n24706,
         p_wishbone_bd_ram_n24707, p_wishbone_bd_ram_n24708,
         p_wishbone_bd_ram_n24709, p_wishbone_bd_ram_n24710,
         p_wishbone_bd_ram_n24711, p_wishbone_bd_ram_n24712,
         p_wishbone_bd_ram_n24713, p_wishbone_bd_ram_n24714,
         p_wishbone_bd_ram_n24715, p_wishbone_bd_ram_n24716,
         p_wishbone_bd_ram_n24717, p_wishbone_bd_ram_n24718,
         p_wishbone_bd_ram_n24719, p_wishbone_bd_ram_n24720,
         p_wishbone_bd_ram_n24721, p_wishbone_bd_ram_n24722,
         p_wishbone_bd_ram_n24723, p_wishbone_bd_ram_n24724,
         p_wishbone_bd_ram_n24725, p_wishbone_bd_ram_n24726,
         p_wishbone_bd_ram_n24727, p_wishbone_bd_ram_n24728,
         p_wishbone_bd_ram_n24729, p_wishbone_bd_ram_n24730,
         p_wishbone_bd_ram_n24731, p_wishbone_bd_ram_n24732,
         p_wishbone_bd_ram_n24733, p_wishbone_bd_ram_n24734,
         p_wishbone_bd_ram_n24735, p_wishbone_bd_ram_n24736,
         p_wishbone_bd_ram_n24737, p_wishbone_bd_ram_n24738,
         p_wishbone_bd_ram_n24739, p_wishbone_bd_ram_n24740,
         p_wishbone_bd_ram_n24741, p_wishbone_bd_ram_n24742,
         p_wishbone_bd_ram_n24743, p_wishbone_bd_ram_n24744,
         p_wishbone_bd_ram_n24745, p_wishbone_bd_ram_n24746,
         p_wishbone_bd_ram_n24747, p_wishbone_bd_ram_n24748,
         p_wishbone_bd_ram_n24749, p_wishbone_bd_ram_n24750,
         p_wishbone_bd_ram_n24751, p_wishbone_bd_ram_n24752,
         p_wishbone_bd_ram_n24753, p_wishbone_bd_ram_n24754,
         p_wishbone_bd_ram_n24755, p_wishbone_bd_ram_n24756,
         p_wishbone_bd_ram_n24757, p_wishbone_bd_ram_n24758,
         p_wishbone_bd_ram_n24759, p_wishbone_bd_ram_n24760,
         p_wishbone_bd_ram_n24761, p_wishbone_bd_ram_n24762,
         p_wishbone_bd_ram_n24763, p_wishbone_bd_ram_n24764,
         p_wishbone_bd_ram_n24765, p_wishbone_bd_ram_n24766,
         p_wishbone_bd_ram_n24767, p_wishbone_bd_ram_n24768,
         p_wishbone_bd_ram_n24769, p_wishbone_bd_ram_n24770,
         p_wishbone_bd_ram_n24771, p_wishbone_bd_ram_n24772,
         p_wishbone_bd_ram_n24773, p_wishbone_bd_ram_n24774,
         p_wishbone_bd_ram_n24775, p_wishbone_bd_ram_n24776,
         p_wishbone_bd_ram_n24777, p_wishbone_bd_ram_n24778,
         p_wishbone_bd_ram_n24779, p_wishbone_bd_ram_n24780,
         p_wishbone_bd_ram_n24781, p_wishbone_bd_ram_n24782,
         p_wishbone_bd_ram_n24783, p_wishbone_bd_ram_n24784,
         p_wishbone_bd_ram_n24785, p_wishbone_bd_ram_n24786,
         p_wishbone_bd_ram_n24787, p_wishbone_bd_ram_n24788,
         p_wishbone_bd_ram_n24789, p_wishbone_bd_ram_n24790,
         p_wishbone_bd_ram_n24791, p_wishbone_bd_ram_n24792,
         p_wishbone_bd_ram_n24793, p_wishbone_bd_ram_n24794,
         p_wishbone_bd_ram_n24795, p_wishbone_bd_ram_n24796,
         p_wishbone_bd_ram_n24797, p_wishbone_bd_ram_n24798,
         p_wishbone_bd_ram_n24799, p_wishbone_bd_ram_n24800,
         p_wishbone_bd_ram_n24801, p_wishbone_bd_ram_n24802,
         p_wishbone_bd_ram_n24803, p_wishbone_bd_ram_n24804,
         p_wishbone_bd_ram_n24805, p_wishbone_bd_ram_n24806,
         p_wishbone_bd_ram_n24807, p_wishbone_bd_ram_n24808,
         p_wishbone_bd_ram_n24809, p_wishbone_bd_ram_n24810,
         p_wishbone_bd_ram_n24811, p_wishbone_bd_ram_n24812,
         p_wishbone_bd_ram_n24813, p_wishbone_bd_ram_n24814,
         p_wishbone_bd_ram_n24815, p_wishbone_bd_ram_n24816,
         p_wishbone_bd_ram_n24817, p_wishbone_bd_ram_n24818,
         p_wishbone_bd_ram_n24819, p_wishbone_bd_ram_n24820,
         p_wishbone_bd_ram_n24821, p_wishbone_bd_ram_n24822,
         p_wishbone_bd_ram_n24823, p_wishbone_bd_ram_n24824,
         p_wishbone_bd_ram_n24825, p_wishbone_bd_ram_n24826,
         p_wishbone_bd_ram_n24827, p_wishbone_bd_ram_n24828,
         p_wishbone_bd_ram_n24829, p_wishbone_bd_ram_n24830,
         p_wishbone_bd_ram_n24831, p_wishbone_bd_ram_n24832,
         p_wishbone_bd_ram_n24833, p_wishbone_bd_ram_n24834,
         p_wishbone_bd_ram_n24835, p_wishbone_bd_ram_n24836,
         p_wishbone_bd_ram_n24837, p_wishbone_bd_ram_n24838,
         p_wishbone_bd_ram_n24839, p_wishbone_bd_ram_n24840,
         p_wishbone_bd_ram_n24841, p_wishbone_bd_ram_n24842,
         p_wishbone_bd_ram_n24843, p_wishbone_bd_ram_n24844,
         p_wishbone_bd_ram_n24845, p_wishbone_bd_ram_n24846,
         p_wishbone_bd_ram_n24847, p_wishbone_bd_ram_n24848,
         p_wishbone_bd_ram_n24849, p_wishbone_bd_ram_n24850,
         p_wishbone_bd_ram_n24851, p_wishbone_bd_ram_n24852,
         p_wishbone_bd_ram_n24853, p_wishbone_bd_ram_n24854,
         p_wishbone_bd_ram_n24855, p_wishbone_bd_ram_n24856,
         p_wishbone_bd_ram_n24857, p_wishbone_bd_ram_n24858,
         p_wishbone_bd_ram_n24859, p_wishbone_bd_ram_n24860,
         p_wishbone_bd_ram_n24861, p_wishbone_bd_ram_n24862,
         p_wishbone_bd_ram_n24863, p_wishbone_bd_ram_n24864,
         p_wishbone_bd_ram_n24865, p_wishbone_bd_ram_n24866,
         p_wishbone_bd_ram_n24867, p_wishbone_bd_ram_n24868,
         p_wishbone_bd_ram_n24869, p_wishbone_bd_ram_n24870,
         p_wishbone_bd_ram_n24871, p_wishbone_bd_ram_n24872,
         p_wishbone_bd_ram_n24873, p_wishbone_bd_ram_n24874,
         p_wishbone_bd_ram_n24875, p_wishbone_bd_ram_n24876,
         p_wishbone_bd_ram_n24877, p_wishbone_bd_ram_n24878,
         p_wishbone_bd_ram_n24879, p_wishbone_bd_ram_n24880,
         p_wishbone_bd_ram_n24881, p_wishbone_bd_ram_n24882,
         p_wishbone_bd_ram_n24883, p_wishbone_bd_ram_n24884,
         p_wishbone_bd_ram_n24885, p_wishbone_bd_ram_n24886,
         p_wishbone_bd_ram_n24887, p_wishbone_bd_ram_n24888,
         p_wishbone_bd_ram_n24889, p_wishbone_bd_ram_n24890,
         p_wishbone_bd_ram_n24891, p_wishbone_bd_ram_n24892,
         p_wishbone_bd_ram_n24893, p_wishbone_bd_ram_n24894,
         p_wishbone_bd_ram_n24895, p_wishbone_bd_ram_n24896,
         p_wishbone_bd_ram_n24897, p_wishbone_bd_ram_n24898,
         p_wishbone_bd_ram_n24899, p_wishbone_bd_ram_n24900,
         p_wishbone_bd_ram_n24901, p_wishbone_bd_ram_n24902,
         p_wishbone_bd_ram_n24903, p_wishbone_bd_ram_n24904,
         p_wishbone_bd_ram_n24905, p_wishbone_bd_ram_n24906,
         p_wishbone_bd_ram_n24907, p_wishbone_bd_ram_n24908,
         p_wishbone_bd_ram_n24909, p_wishbone_bd_ram_n24910,
         p_wishbone_bd_ram_n24911, p_wishbone_bd_ram_n24912,
         p_wishbone_bd_ram_n24913, p_wishbone_bd_ram_n24914,
         p_wishbone_bd_ram_n24915, p_wishbone_bd_ram_n24916,
         p_wishbone_bd_ram_n24917, p_wishbone_bd_ram_n24918,
         p_wishbone_bd_ram_n24919, p_wishbone_bd_ram_n24920,
         p_wishbone_bd_ram_n24921, p_wishbone_bd_ram_n24922,
         p_wishbone_bd_ram_n24923, p_wishbone_bd_ram_n24924,
         p_wishbone_bd_ram_n24925, p_wishbone_bd_ram_n24926,
         p_wishbone_bd_ram_n24927, p_wishbone_bd_ram_n24928,
         p_wishbone_bd_ram_n24929, p_wishbone_bd_ram_n24930,
         p_wishbone_bd_ram_n24931, p_wishbone_bd_ram_n24932,
         p_wishbone_bd_ram_n24933, p_wishbone_bd_ram_n24934,
         p_wishbone_bd_ram_n24935, p_wishbone_bd_ram_n24936,
         p_wishbone_bd_ram_n24937, p_wishbone_bd_ram_n24938,
         p_wishbone_bd_ram_n24939, p_wishbone_bd_ram_n24940,
         p_wishbone_bd_ram_n24941, p_wishbone_bd_ram_n24942,
         p_wishbone_bd_ram_n24943, p_wishbone_bd_ram_n24944,
         p_wishbone_bd_ram_n24945, p_wishbone_bd_ram_n24946,
         p_wishbone_bd_ram_n24947, p_wishbone_bd_ram_n24948,
         p_wishbone_bd_ram_n24949, p_wishbone_bd_ram_n24950,
         p_wishbone_bd_ram_n24951, p_wishbone_bd_ram_n24952,
         p_wishbone_bd_ram_n24953, p_wishbone_bd_ram_n24954,
         p_wishbone_bd_ram_n24955, p_wishbone_bd_ram_n24956,
         p_wishbone_bd_ram_n24957, p_wishbone_bd_ram_n24958,
         p_wishbone_bd_ram_n24959, p_wishbone_bd_ram_n24960,
         p_wishbone_bd_ram_n24961, p_wishbone_bd_ram_n24962,
         p_wishbone_bd_ram_n24963, p_wishbone_bd_ram_n24964,
         p_wishbone_bd_ram_n24965, p_wishbone_bd_ram_n24966,
         p_wishbone_bd_ram_n24967, p_wishbone_bd_ram_n24968,
         p_wishbone_bd_ram_n24969, p_wishbone_bd_ram_n24970,
         p_wishbone_bd_ram_n24971, p_wishbone_bd_ram_n24972,
         p_wishbone_bd_ram_n24973, p_wishbone_bd_ram_n24974,
         p_wishbone_bd_ram_n24975, p_wishbone_bd_ram_n24976,
         p_wishbone_bd_ram_n24977, p_wishbone_bd_ram_n24978,
         p_wishbone_bd_ram_n24979, p_wishbone_bd_ram_n24980,
         p_wishbone_bd_ram_n24981, p_wishbone_bd_ram_n24982,
         p_wishbone_bd_ram_n24983, p_wishbone_bd_ram_n24984,
         p_wishbone_bd_ram_n24985, p_wishbone_bd_ram_n24986,
         p_wishbone_bd_ram_n24987, p_wishbone_bd_ram_n24988,
         p_wishbone_bd_ram_n24989, p_wishbone_bd_ram_n24990,
         p_wishbone_bd_ram_n24991, p_wishbone_bd_ram_n24992,
         p_wishbone_bd_ram_n24993, p_wishbone_bd_ram_n24994,
         p_wishbone_bd_ram_n24995, p_wishbone_bd_ram_n24996,
         p_wishbone_bd_ram_n24997, p_wishbone_bd_ram_n24998,
         p_wishbone_bd_ram_n24999, p_wishbone_bd_ram_n25000,
         p_wishbone_bd_ram_n25001, p_wishbone_bd_ram_n25002,
         p_wishbone_bd_ram_n25003, p_wishbone_bd_ram_n25004,
         p_wishbone_bd_ram_n25005, p_wishbone_bd_ram_n25006,
         p_wishbone_bd_ram_n25007, p_wishbone_bd_ram_n25008,
         p_wishbone_bd_ram_n25009, p_wishbone_bd_ram_n25010,
         p_wishbone_bd_ram_n25011, p_wishbone_bd_ram_n25012,
         p_wishbone_bd_ram_n25013, p_wishbone_bd_ram_n25014,
         p_wishbone_bd_ram_n25015, p_wishbone_bd_ram_n25016,
         p_wishbone_bd_ram_n25017, p_wishbone_bd_ram_n25018,
         p_wishbone_bd_ram_n25019, p_wishbone_bd_ram_n25020,
         p_wishbone_bd_ram_n25021, p_wishbone_bd_ram_n25022,
         p_wishbone_bd_ram_n25023, p_wishbone_bd_ram_n25024,
         p_wishbone_bd_ram_n25025, p_wishbone_bd_ram_n25026,
         p_wishbone_bd_ram_n25027, p_wishbone_bd_ram_n25028,
         p_wishbone_bd_ram_n25029, p_wishbone_bd_ram_n25030,
         p_wishbone_bd_ram_n25031, p_wishbone_bd_ram_n25032,
         p_wishbone_bd_ram_n25033, p_wishbone_bd_ram_n25034,
         p_wishbone_bd_ram_n25035, p_wishbone_bd_ram_n25036,
         p_wishbone_bd_ram_n25037, p_wishbone_bd_ram_n25038,
         p_wishbone_bd_ram_n25039, p_wishbone_bd_ram_n25040,
         p_wishbone_bd_ram_n25041, p_wishbone_bd_ram_n25042,
         p_wishbone_bd_ram_n25043, p_wishbone_bd_ram_n25044,
         p_wishbone_bd_ram_n25045, p_wishbone_bd_ram_n25046,
         p_wishbone_bd_ram_n25047, p_wishbone_bd_ram_n25048,
         p_wishbone_bd_ram_n25049, p_wishbone_bd_ram_n25050,
         p_wishbone_bd_ram_n25051, p_wishbone_bd_ram_n25052,
         p_wishbone_bd_ram_n25053, p_wishbone_bd_ram_n25054,
         p_wishbone_bd_ram_n25055, p_wishbone_bd_ram_n25056,
         p_wishbone_bd_ram_n25057, p_wishbone_bd_ram_n25058,
         p_wishbone_bd_ram_n25059, p_wishbone_bd_ram_n25060,
         p_wishbone_bd_ram_n25061, p_wishbone_bd_ram_n25062,
         p_wishbone_bd_ram_n25063, p_wishbone_bd_ram_n25064,
         p_wishbone_bd_ram_n25065, p_wishbone_bd_ram_n25066,
         p_wishbone_bd_ram_n25067, p_wishbone_bd_ram_n25068,
         p_wishbone_bd_ram_n25069, p_wishbone_bd_ram_n25070,
         p_wishbone_bd_ram_n25071, p_wishbone_bd_ram_n25072,
         p_wishbone_bd_ram_n25073, p_wishbone_bd_ram_n25074,
         p_wishbone_bd_ram_n25075, p_wishbone_bd_ram_n25076,
         p_wishbone_bd_ram_n25077, p_wishbone_bd_ram_n25078,
         p_wishbone_bd_ram_n25079, p_wishbone_bd_ram_n25080,
         p_wishbone_bd_ram_n25081, p_wishbone_bd_ram_n25082,
         p_wishbone_bd_ram_n25083, p_wishbone_bd_ram_n25084,
         p_wishbone_bd_ram_n25085, p_wishbone_bd_ram_n25086,
         p_wishbone_bd_ram_n25087, p_wishbone_bd_ram_n25088,
         p_wishbone_bd_ram_n25089, p_wishbone_bd_ram_n25090,
         p_wishbone_bd_ram_n25091, p_wishbone_bd_ram_n25092,
         p_wishbone_bd_ram_n25093, p_wishbone_bd_ram_n25094,
         p_wishbone_bd_ram_n25095, p_wishbone_bd_ram_n25096,
         p_wishbone_bd_ram_n25097, p_wishbone_bd_ram_n25098,
         p_wishbone_bd_ram_n25099, p_wishbone_bd_ram_n25100,
         p_wishbone_bd_ram_n25101, p_wishbone_bd_ram_n25102,
         p_wishbone_bd_ram_n25103, p_wishbone_bd_ram_n25104,
         p_wishbone_bd_ram_n25105, p_wishbone_bd_ram_n25106,
         p_wishbone_bd_ram_n25107, p_wishbone_bd_ram_n25108,
         p_wishbone_bd_ram_n25109, p_wishbone_bd_ram_n25110,
         p_wishbone_bd_ram_n25111, p_wishbone_bd_ram_n25112,
         p_wishbone_bd_ram_n25113, p_wishbone_bd_ram_n25114,
         p_wishbone_bd_ram_n25115, p_wishbone_bd_ram_n25116,
         p_wishbone_bd_ram_n25117, p_wishbone_bd_ram_n25118,
         p_wishbone_bd_ram_n25119, p_wishbone_bd_ram_n25120,
         p_wishbone_bd_ram_n25121, p_wishbone_bd_ram_n25122,
         p_wishbone_bd_ram_n25123, p_wishbone_bd_ram_n25124,
         p_wishbone_bd_ram_n25125, p_wishbone_bd_ram_n25126,
         p_wishbone_bd_ram_n25127, p_wishbone_bd_ram_n25128,
         p_wishbone_bd_ram_n25129, p_wishbone_bd_ram_n25130,
         p_wishbone_bd_ram_n25131, p_wishbone_bd_ram_n25132,
         p_wishbone_bd_ram_n25133, p_wishbone_bd_ram_n25134,
         p_wishbone_bd_ram_n25135, p_wishbone_bd_ram_n25136,
         p_wishbone_bd_ram_n25137, p_wishbone_bd_ram_n25138,
         p_wishbone_bd_ram_n25139, p_wishbone_bd_ram_n25140,
         p_wishbone_bd_ram_n25141, p_wishbone_bd_ram_n25142,
         p_wishbone_bd_ram_n25143, p_wishbone_bd_ram_n25144,
         p_wishbone_bd_ram_n25145, p_wishbone_bd_ram_n25146,
         p_wishbone_bd_ram_n25147, p_wishbone_bd_ram_n25148,
         p_wishbone_bd_ram_n25149, p_wishbone_bd_ram_n25150,
         p_wishbone_bd_ram_n25151, p_wishbone_bd_ram_n25152,
         p_wishbone_bd_ram_n25153, p_wishbone_bd_ram_n25154,
         p_wishbone_bd_ram_n25155, p_wishbone_bd_ram_n25156,
         p_wishbone_bd_ram_n25157, p_wishbone_bd_ram_n25158,
         p_wishbone_bd_ram_n25159, p_wishbone_bd_ram_n25160,
         p_wishbone_bd_ram_n25161, p_wishbone_bd_ram_n25162,
         p_wishbone_bd_ram_n25163, p_wishbone_bd_ram_n25164,
         p_wishbone_bd_ram_n25165, p_wishbone_bd_ram_n25166,
         p_wishbone_bd_ram_n25167, p_wishbone_bd_ram_n25168,
         p_wishbone_bd_ram_n25169, p_wishbone_bd_ram_n25170,
         p_wishbone_bd_ram_n25171, p_wishbone_bd_ram_n25172,
         p_wishbone_bd_ram_n25173, p_wishbone_bd_ram_n25174,
         p_wishbone_bd_ram_n25175, p_wishbone_bd_ram_n25176,
         p_wishbone_bd_ram_n25177, p_wishbone_bd_ram_n25178,
         p_wishbone_bd_ram_n25179, p_wishbone_bd_ram_n25180,
         p_wishbone_bd_ram_n25181, p_wishbone_bd_ram_n25182,
         p_wishbone_bd_ram_n25183, p_wishbone_bd_ram_n25184,
         p_wishbone_bd_ram_n25185, p_wishbone_bd_ram_n25186,
         p_wishbone_bd_ram_n25187, p_wishbone_bd_ram_n25188,
         p_wishbone_bd_ram_n25189, p_wishbone_bd_ram_n25190,
         p_wishbone_bd_ram_n25191, p_wishbone_bd_ram_n25192,
         p_wishbone_bd_ram_n25193, p_wishbone_bd_ram_n25194,
         p_wishbone_bd_ram_n25195, p_wishbone_bd_ram_n25196,
         p_wishbone_bd_ram_n25197, p_wishbone_bd_ram_n25198,
         p_wishbone_bd_ram_n25199, p_wishbone_bd_ram_n25200,
         p_wishbone_bd_ram_n25201, p_wishbone_bd_ram_n25202,
         p_wishbone_bd_ram_n25203, p_wishbone_bd_ram_n25204,
         p_wishbone_bd_ram_n25205, p_wishbone_bd_ram_n25206,
         p_wishbone_bd_ram_n25207, p_wishbone_bd_ram_n25208,
         p_wishbone_bd_ram_n25209, p_wishbone_bd_ram_n25210,
         p_wishbone_bd_ram_n25211, p_wishbone_bd_ram_n25212,
         p_wishbone_bd_ram_n25213, p_wishbone_bd_ram_n25214,
         p_wishbone_bd_ram_n25215, p_wishbone_bd_ram_n25216,
         p_wishbone_bd_ram_n25217, p_wishbone_bd_ram_n25218,
         p_wishbone_bd_ram_n25219, p_wishbone_bd_ram_n25220,
         p_wishbone_bd_ram_n25221, p_wishbone_bd_ram_n25222,
         p_wishbone_bd_ram_n25223, p_wishbone_bd_ram_n25224,
         p_wishbone_bd_ram_n25225, p_wishbone_bd_ram_n25226,
         p_wishbone_bd_ram_n25227, p_wishbone_bd_ram_n25228,
         p_wishbone_bd_ram_n25229, p_wishbone_bd_ram_n25230,
         p_wishbone_bd_ram_n25231, p_wishbone_bd_ram_n25232,
         p_wishbone_bd_ram_n25233, p_wishbone_bd_ram_n25234,
         p_wishbone_bd_ram_n25235, p_wishbone_bd_ram_n25236,
         p_wishbone_bd_ram_n25237, p_wishbone_bd_ram_n25238,
         p_wishbone_bd_ram_n25239, p_wishbone_bd_ram_n25240,
         p_wishbone_bd_ram_n25241, p_wishbone_bd_ram_n25242,
         p_wishbone_bd_ram_n25243, p_wishbone_bd_ram_n25244,
         p_wishbone_bd_ram_n25245, p_wishbone_bd_ram_n25246,
         p_wishbone_bd_ram_n25247, p_wishbone_bd_ram_n25248,
         p_wishbone_bd_ram_n25249, p_wishbone_bd_ram_n25250,
         p_wishbone_bd_ram_n25251, p_wishbone_bd_ram_n25252,
         p_wishbone_bd_ram_n25253, p_wishbone_bd_ram_n25254,
         p_wishbone_bd_ram_n25255, p_wishbone_bd_ram_n25256,
         p_wishbone_bd_ram_n25257, p_wishbone_bd_ram_n25258,
         p_wishbone_bd_ram_n25259, p_wishbone_bd_ram_n25260,
         p_wishbone_bd_ram_n25261, p_wishbone_bd_ram_n25262,
         p_wishbone_bd_ram_n25263, p_wishbone_bd_ram_n25264,
         p_wishbone_bd_ram_n25265, p_wishbone_bd_ram_n25266,
         p_wishbone_bd_ram_n25267, p_wishbone_bd_ram_n25268,
         p_wishbone_bd_ram_n25269, p_wishbone_bd_ram_n25270,
         p_wishbone_bd_ram_n25271, p_wishbone_bd_ram_n25272,
         p_wishbone_bd_ram_n25273, p_wishbone_bd_ram_n25274,
         p_wishbone_bd_ram_n25275, p_wishbone_bd_ram_n25276,
         p_wishbone_bd_ram_n25277, p_wishbone_bd_ram_n25278,
         p_wishbone_bd_ram_n25279, p_wishbone_bd_ram_n25280,
         p_wishbone_bd_ram_n25281, p_wishbone_bd_ram_n25282,
         p_wishbone_bd_ram_n25283, p_wishbone_bd_ram_n25284,
         p_wishbone_bd_ram_n25285, p_wishbone_bd_ram_n25286,
         p_wishbone_bd_ram_n25287, p_wishbone_bd_ram_n25288,
         p_wishbone_bd_ram_n25289, p_wishbone_bd_ram_n25290,
         p_wishbone_bd_ram_n25291, p_wishbone_bd_ram_n25292,
         p_wishbone_bd_ram_n25293, p_wishbone_bd_ram_n25294,
         p_wishbone_bd_ram_n25295, p_wishbone_bd_ram_n25296,
         p_wishbone_bd_ram_n25297, p_wishbone_bd_ram_n25298,
         p_wishbone_bd_ram_n25299, p_wishbone_bd_ram_n25300,
         p_wishbone_bd_ram_n25301, p_wishbone_bd_ram_n25302,
         p_wishbone_bd_ram_n25303, p_wishbone_bd_ram_n25304,
         p_wishbone_bd_ram_n25305, p_wishbone_bd_ram_n25306,
         p_wishbone_bd_ram_n25307, p_wishbone_bd_ram_n25308,
         p_wishbone_bd_ram_n25309, p_wishbone_bd_ram_n25310,
         p_wishbone_bd_ram_n25311, p_wishbone_bd_ram_n25312,
         p_wishbone_bd_ram_n25313, p_wishbone_bd_ram_n25314,
         p_wishbone_bd_ram_n25315, p_wishbone_bd_ram_n25316,
         p_wishbone_bd_ram_n25317, p_wishbone_bd_ram_n25318,
         p_wishbone_bd_ram_n25319, p_wishbone_bd_ram_n25320,
         p_wishbone_bd_ram_n25321, p_wishbone_bd_ram_n25322,
         p_wishbone_bd_ram_n25323, p_wishbone_bd_ram_n25324,
         p_wishbone_bd_ram_n25325, p_wishbone_bd_ram_n25326,
         p_wishbone_bd_ram_n25327, p_wishbone_bd_ram_n25328,
         p_wishbone_bd_ram_n25329, p_wishbone_bd_ram_n25330,
         p_wishbone_bd_ram_n25331, p_wishbone_bd_ram_n25332,
         p_wishbone_bd_ram_n25333, p_wishbone_bd_ram_n25334,
         p_wishbone_bd_ram_n25335, p_wishbone_bd_ram_n25336,
         p_wishbone_bd_ram_n25337, p_wishbone_bd_ram_n25338,
         p_wishbone_bd_ram_n25339, p_wishbone_bd_ram_n25340,
         p_wishbone_bd_ram_n25341, p_wishbone_bd_ram_n25342,
         p_wishbone_bd_ram_n25343, p_wishbone_bd_ram_n25344,
         p_wishbone_bd_ram_n25345, p_wishbone_bd_ram_n25346,
         p_wishbone_bd_ram_n25347, p_wishbone_bd_ram_n25348,
         p_wishbone_bd_ram_n25349, p_wishbone_bd_ram_n25350,
         p_wishbone_bd_ram_n25351, p_wishbone_bd_ram_n25352,
         p_wishbone_bd_ram_n25353, p_wishbone_bd_ram_n25354,
         p_wishbone_bd_ram_n25355, p_wishbone_bd_ram_n25356,
         p_wishbone_bd_ram_n25357, p_wishbone_bd_ram_n25358,
         p_wishbone_bd_ram_n25359, p_wishbone_bd_ram_n25360,
         p_wishbone_bd_ram_n25361, p_wishbone_bd_ram_n25362,
         p_wishbone_bd_ram_n25363, p_wishbone_bd_ram_n25364,
         p_wishbone_bd_ram_n25365, p_wishbone_bd_ram_n25366,
         p_wishbone_bd_ram_n25367, p_wishbone_bd_ram_n25368,
         p_wishbone_bd_ram_n25369, p_wishbone_bd_ram_n25370,
         p_wishbone_bd_ram_n25371, p_wishbone_bd_ram_n25372,
         p_wishbone_bd_ram_n25373, p_wishbone_bd_ram_n25374,
         p_wishbone_bd_ram_n25375, p_wishbone_bd_ram_n25376,
         p_wishbone_bd_ram_n25377, p_wishbone_bd_ram_n25378,
         p_wishbone_bd_ram_n25379, p_wishbone_bd_ram_n25380,
         p_wishbone_bd_ram_n25381, p_wishbone_bd_ram_n25382,
         p_wishbone_bd_ram_n25383, p_wishbone_bd_ram_n25384,
         p_wishbone_bd_ram_n25385, p_wishbone_bd_ram_n25386,
         p_wishbone_bd_ram_n25387, p_wishbone_bd_ram_n25388,
         p_wishbone_bd_ram_n25389, p_wishbone_bd_ram_n25390,
         p_wishbone_bd_ram_n25391, p_wishbone_bd_ram_n25392,
         p_wishbone_bd_ram_n25393, p_wishbone_bd_ram_n25394,
         p_wishbone_bd_ram_n25395, p_wishbone_bd_ram_n25396,
         p_wishbone_bd_ram_n25397, p_wishbone_bd_ram_n25398,
         p_wishbone_bd_ram_n25399, p_wishbone_bd_ram_n25400,
         p_wishbone_bd_ram_n25401, p_wishbone_bd_ram_n25402,
         p_wishbone_bd_ram_n25403, p_wishbone_bd_ram_n25404,
         p_wishbone_bd_ram_n25405, p_wishbone_bd_ram_n25406,
         p_wishbone_bd_ram_n25407, p_wishbone_bd_ram_n25408,
         p_wishbone_bd_ram_n25409, p_wishbone_bd_ram_n25410,
         p_wishbone_bd_ram_n25411, p_wishbone_bd_ram_n25412,
         p_wishbone_bd_ram_n25413, p_wishbone_bd_ram_n25414,
         p_wishbone_bd_ram_n25415, p_wishbone_bd_ram_n25416,
         p_wishbone_bd_ram_n25417, p_wishbone_bd_ram_n25418,
         p_wishbone_bd_ram_n25419, p_wishbone_bd_ram_n25420,
         p_wishbone_bd_ram_n25421, p_wishbone_bd_ram_n25422,
         p_wishbone_bd_ram_n25423, p_wishbone_bd_ram_n25424,
         p_wishbone_bd_ram_n25425, p_wishbone_bd_ram_n25426,
         p_wishbone_bd_ram_n25427, p_wishbone_bd_ram_n25428,
         p_wishbone_bd_ram_n25429, p_wishbone_bd_ram_n25430,
         p_wishbone_bd_ram_n25431, p_wishbone_bd_ram_n25432,
         p_wishbone_bd_ram_n25433, p_wishbone_bd_ram_n25434,
         p_wishbone_bd_ram_n25435, p_wishbone_bd_ram_n25436,
         p_wishbone_bd_ram_n25437, p_wishbone_bd_ram_n25438,
         p_wishbone_bd_ram_n25439, p_wishbone_bd_ram_n25440,
         p_wishbone_bd_ram_n25441, p_wishbone_bd_ram_n25442,
         p_wishbone_bd_ram_n25443, p_wishbone_bd_ram_n25444,
         p_wishbone_bd_ram_n25445, p_wishbone_bd_ram_n25446,
         p_wishbone_bd_ram_n25447, p_wishbone_bd_ram_n25448,
         p_wishbone_bd_ram_n25449, p_wishbone_bd_ram_n25450,
         p_wishbone_bd_ram_n25451, p_wishbone_bd_ram_n25452,
         p_wishbone_bd_ram_n25453, p_wishbone_bd_ram_n25454,
         p_wishbone_bd_ram_n25455, p_wishbone_bd_ram_n25456,
         p_wishbone_bd_ram_n25457, p_wishbone_bd_ram_n25458,
         p_wishbone_bd_ram_n25459, p_wishbone_bd_ram_n25460,
         p_wishbone_bd_ram_n25461, p_wishbone_bd_ram_n25462,
         p_wishbone_bd_ram_n25463, p_wishbone_bd_ram_n25464,
         p_wishbone_bd_ram_n25465, p_wishbone_bd_ram_n25466,
         p_wishbone_bd_ram_n25467, p_wishbone_bd_ram_n25468,
         p_wishbone_bd_ram_n25469, p_wishbone_bd_ram_n25470,
         p_wishbone_bd_ram_n25471, p_wishbone_bd_ram_n25472,
         p_wishbone_bd_ram_n25473, p_wishbone_bd_ram_n25474,
         p_wishbone_bd_ram_n25475, p_wishbone_bd_ram_n25476,
         p_wishbone_bd_ram_n25477, p_wishbone_bd_ram_n25478,
         p_wishbone_bd_ram_n25479, p_wishbone_bd_ram_n25480,
         p_wishbone_bd_ram_n25481, p_wishbone_bd_ram_n25482,
         p_wishbone_bd_ram_n25483, p_wishbone_bd_ram_n25484,
         p_wishbone_bd_ram_n25485, p_wishbone_bd_ram_n25486,
         p_wishbone_bd_ram_n25487, p_wishbone_bd_ram_n25488,
         p_wishbone_bd_ram_n25489, p_wishbone_bd_ram_n25490,
         p_wishbone_bd_ram_n25491, p_wishbone_bd_ram_n25492,
         p_wishbone_bd_ram_n25493, p_wishbone_bd_ram_n25494,
         p_wishbone_bd_ram_n25495, p_wishbone_bd_ram_n25496,
         p_wishbone_bd_ram_n25497, p_wishbone_bd_ram_n25498,
         p_wishbone_bd_ram_n25499, p_wishbone_bd_ram_n25500,
         p_wishbone_bd_ram_n25501, p_wishbone_bd_ram_n25502,
         p_wishbone_bd_ram_n25503, p_wishbone_bd_ram_n25504,
         p_wishbone_bd_ram_n25505, p_wishbone_bd_ram_n25506,
         p_wishbone_bd_ram_n25507, p_wishbone_bd_ram_n25508,
         p_wishbone_bd_ram_n25509, p_wishbone_bd_ram_n25510,
         p_wishbone_bd_ram_n25511, p_wishbone_bd_ram_n25512,
         p_wishbone_bd_ram_n25513, p_wishbone_bd_ram_n25514,
         p_wishbone_bd_ram_n25515, p_wishbone_bd_ram_n25516,
         p_wishbone_bd_ram_n25517, p_wishbone_bd_ram_n25518,
         p_wishbone_bd_ram_n25519, p_wishbone_bd_ram_n25520,
         p_wishbone_bd_ram_n25521, p_wishbone_bd_ram_n25522,
         p_wishbone_bd_ram_n25523, p_wishbone_bd_ram_n25524,
         p_wishbone_bd_ram_n25525, p_wishbone_bd_ram_n25526,
         p_wishbone_bd_ram_n25527, p_wishbone_bd_ram_n25528,
         p_wishbone_bd_ram_n25529, p_wishbone_bd_ram_n25530,
         p_wishbone_bd_ram_n25531, p_wishbone_bd_ram_n25532,
         p_wishbone_bd_ram_n25533, p_wishbone_bd_ram_n25534,
         p_wishbone_bd_ram_n25535, p_wishbone_bd_ram_n25536,
         p_wishbone_bd_ram_n25537, p_wishbone_bd_ram_n25538,
         p_wishbone_bd_ram_n25539, p_wishbone_bd_ram_n25540,
         p_wishbone_bd_ram_n25541, p_wishbone_bd_ram_n25542,
         p_wishbone_bd_ram_n25543, p_wishbone_bd_ram_n25544,
         p_wishbone_bd_ram_n25545, p_wishbone_bd_ram_n25546,
         p_wishbone_bd_ram_n25547, p_wishbone_bd_ram_n25548,
         p_wishbone_bd_ram_n25549, p_wishbone_bd_ram_n25550,
         p_wishbone_bd_ram_n25551, p_wishbone_bd_ram_n25552,
         p_wishbone_bd_ram_n25553, p_wishbone_bd_ram_n25554,
         p_wishbone_bd_ram_n25555, p_wishbone_bd_ram_n25556,
         p_wishbone_bd_ram_n25557, p_wishbone_bd_ram_n25558,
         p_wishbone_bd_ram_n25559, p_wishbone_bd_ram_n25560,
         p_wishbone_bd_ram_n25561, p_wishbone_bd_ram_n25562,
         p_wishbone_bd_ram_n25563, p_wishbone_bd_ram_n25564,
         p_wishbone_bd_ram_n25565, p_wishbone_bd_ram_n25566,
         p_wishbone_bd_ram_n25567, p_wishbone_bd_ram_n25568,
         p_wishbone_bd_ram_n25569, p_wishbone_bd_ram_n25570,
         p_wishbone_bd_ram_n25571, p_wishbone_bd_ram_n25572,
         p_wishbone_bd_ram_n25573, p_wishbone_bd_ram_n25574,
         p_wishbone_bd_ram_n25575, p_wishbone_bd_ram_n25576,
         p_wishbone_bd_ram_n25577, p_wishbone_bd_ram_n25578,
         p_wishbone_bd_ram_n25579, p_wishbone_bd_ram_n25580,
         p_wishbone_bd_ram_n25581, p_wishbone_bd_ram_n25582,
         p_wishbone_bd_ram_n25583, p_wishbone_bd_ram_n25584,
         p_wishbone_bd_ram_n25585, p_wishbone_bd_ram_n25586,
         p_wishbone_bd_ram_n25587, p_wishbone_bd_ram_n25588,
         p_wishbone_bd_ram_n25589, p_wishbone_bd_ram_n25590,
         p_wishbone_bd_ram_n25591, p_wishbone_bd_ram_n25592,
         p_wishbone_bd_ram_n25593, p_wishbone_bd_ram_n25594,
         p_wishbone_bd_ram_n25595, p_wishbone_bd_ram_n25596,
         p_wishbone_bd_ram_n25597, p_wishbone_bd_ram_n25598,
         p_wishbone_bd_ram_n25599, p_wishbone_bd_ram_n25600,
         p_wishbone_bd_ram_n25601, p_wishbone_bd_ram_n25602,
         p_wishbone_bd_ram_n25603, p_wishbone_bd_ram_n25604,
         p_wishbone_bd_ram_n25605, p_wishbone_bd_ram_n25606,
         p_wishbone_bd_ram_n25607, p_wishbone_bd_ram_n25608,
         p_wishbone_bd_ram_n25609, p_wishbone_bd_ram_n25610,
         p_wishbone_bd_ram_n25611, p_wishbone_bd_ram_n25612,
         p_wishbone_bd_ram_n25613, p_wishbone_bd_ram_n25614,
         p_wishbone_bd_ram_n25615, p_wishbone_bd_ram_n25616,
         p_wishbone_bd_ram_n25617, p_wishbone_bd_ram_n25618,
         p_wishbone_bd_ram_n25619, p_wishbone_bd_ram_n25620,
         p_wishbone_bd_ram_n25621, p_wishbone_bd_ram_n25622,
         p_wishbone_bd_ram_n25623, p_wishbone_bd_ram_n25624,
         p_wishbone_bd_ram_n25625, p_wishbone_bd_ram_n25626,
         p_wishbone_bd_ram_n25627, p_wishbone_bd_ram_n25628,
         p_wishbone_bd_ram_n25629, p_wishbone_bd_ram_n25630,
         p_wishbone_bd_ram_n25631, p_wishbone_bd_ram_n25632,
         p_wishbone_bd_ram_n25633, p_wishbone_bd_ram_n25634,
         p_wishbone_bd_ram_n25635, p_wishbone_bd_ram_n25636,
         p_wishbone_bd_ram_n25637, p_wishbone_bd_ram_n25638,
         p_wishbone_bd_ram_n25639, p_wishbone_bd_ram_n25640,
         p_wishbone_bd_ram_n25641, p_wishbone_bd_ram_n25642,
         p_wishbone_bd_ram_n25643, p_wishbone_bd_ram_n25644,
         p_wishbone_bd_ram_n25645, p_wishbone_bd_ram_n25646,
         p_wishbone_bd_ram_n25647, p_wishbone_bd_ram_n25648,
         p_wishbone_bd_ram_n25649, p_wishbone_bd_ram_n25650,
         p_wishbone_bd_ram_n25651, p_wishbone_bd_ram_n25652,
         p_wishbone_bd_ram_n25653, p_wishbone_bd_ram_n25654,
         p_wishbone_bd_ram_n25655, p_wishbone_bd_ram_n25656,
         p_wishbone_bd_ram_n25657, p_wishbone_bd_ram_n25658,
         p_wishbone_bd_ram_n25659, p_wishbone_bd_ram_n25660,
         p_wishbone_bd_ram_n25661, p_wishbone_bd_ram_n25662,
         p_wishbone_bd_ram_n25663, p_wishbone_bd_ram_n25664,
         p_wishbone_bd_ram_n25665, p_wishbone_bd_ram_n25666,
         p_wishbone_bd_ram_n25667, p_wishbone_bd_ram_n25668,
         p_wishbone_bd_ram_n25669, p_wishbone_bd_ram_n25670,
         p_wishbone_bd_ram_n25671, p_wishbone_bd_ram_n25672,
         p_wishbone_bd_ram_n25673, p_wishbone_bd_ram_n25674,
         p_wishbone_bd_ram_n25675, p_wishbone_bd_ram_n25676,
         p_wishbone_bd_ram_n25677, p_wishbone_bd_ram_n25678,
         p_wishbone_bd_ram_n25679, p_wishbone_bd_ram_n25680,
         p_wishbone_bd_ram_n25681, p_wishbone_bd_ram_n25682,
         p_wishbone_bd_ram_n25683, p_wishbone_bd_ram_n25684,
         p_wishbone_bd_ram_n25685, p_wishbone_bd_ram_n25686,
         p_wishbone_bd_ram_n25687, p_wishbone_bd_ram_n25688,
         p_wishbone_bd_ram_n25689, p_wishbone_bd_ram_n25690,
         p_wishbone_bd_ram_n25691, p_wishbone_bd_ram_n25692,
         p_wishbone_bd_ram_n25693, p_wishbone_bd_ram_n25694,
         p_wishbone_bd_ram_n25695, p_wishbone_bd_ram_n25696,
         p_wishbone_bd_ram_n25697, p_wishbone_bd_ram_n25698,
         p_wishbone_bd_ram_n25699, p_wishbone_bd_ram_n25700,
         p_wishbone_bd_ram_n25701, p_wishbone_bd_ram_n25702,
         p_wishbone_bd_ram_n25703, p_wishbone_bd_ram_n25704,
         p_wishbone_bd_ram_n25705, p_wishbone_bd_ram_n25706,
         p_wishbone_bd_ram_n25707, p_wishbone_bd_ram_n25708,
         p_wishbone_bd_ram_n25709, p_wishbone_bd_ram_n25710,
         p_wishbone_bd_ram_n25711, p_wishbone_bd_ram_n25712,
         p_wishbone_bd_ram_n25713, p_wishbone_bd_ram_n25714,
         p_wishbone_bd_ram_n25715, p_wishbone_bd_ram_n25716,
         p_wishbone_bd_ram_n25717, p_wishbone_bd_ram_n25718,
         p_wishbone_bd_ram_n25719, p_wishbone_bd_ram_n25720,
         p_wishbone_bd_ram_n25721, p_wishbone_bd_ram_n25722,
         p_wishbone_bd_ram_n25723, p_wishbone_bd_ram_n25724,
         p_wishbone_bd_ram_n25725, p_wishbone_bd_ram_n25726,
         p_wishbone_bd_ram_n25727, p_wishbone_bd_ram_n25728,
         p_wishbone_bd_ram_n25729, p_wishbone_bd_ram_n25730,
         p_wishbone_bd_ram_n25731, p_wishbone_bd_ram_n25732,
         p_wishbone_bd_ram_n25733, p_wishbone_bd_ram_n25734,
         p_wishbone_bd_ram_n25735, p_wishbone_bd_ram_n25736,
         p_wishbone_bd_ram_n25737, p_wishbone_bd_ram_n25738,
         p_wishbone_bd_ram_n25739, p_wishbone_bd_ram_n25740,
         p_wishbone_bd_ram_n25741, p_wishbone_bd_ram_n25742,
         p_wishbone_bd_ram_n25743, p_wishbone_bd_ram_n25744,
         p_wishbone_bd_ram_n25745, p_wishbone_bd_ram_n25746,
         p_wishbone_bd_ram_n25747, p_wishbone_bd_ram_n25748,
         p_wishbone_bd_ram_n25749, p_wishbone_bd_ram_n25750,
         p_wishbone_bd_ram_n25751, p_wishbone_bd_ram_n25752,
         p_wishbone_bd_ram_n25753, p_wishbone_bd_ram_n25754,
         p_wishbone_bd_ram_n25755, p_wishbone_bd_ram_n25756,
         p_wishbone_bd_ram_n25757, p_wishbone_bd_ram_n25758,
         p_wishbone_bd_ram_n25759, p_wishbone_bd_ram_n25760,
         p_wishbone_bd_ram_n25761, p_wishbone_bd_ram_n25762,
         p_wishbone_bd_ram_n25763, p_wishbone_bd_ram_n25764,
         p_wishbone_bd_ram_n25765, p_wishbone_bd_ram_n25766,
         p_wishbone_bd_ram_n25767, p_wishbone_bd_ram_n25768,
         p_wishbone_bd_ram_n25769, p_wishbone_bd_ram_n25770,
         p_wishbone_bd_ram_n25771, p_wishbone_bd_ram_n25772,
         p_wishbone_bd_ram_n25773, p_wishbone_bd_ram_n25774,
         p_wishbone_bd_ram_n25775, p_wishbone_bd_ram_n25776,
         p_wishbone_bd_ram_n25777, p_wishbone_bd_ram_n25778,
         p_wishbone_bd_ram_n25779, p_wishbone_bd_ram_n25780,
         p_wishbone_bd_ram_n25781, p_wishbone_bd_ram_n25782,
         p_wishbone_bd_ram_n25783, p_wishbone_bd_ram_n25784,
         p_wishbone_bd_ram_n25785, p_wishbone_bd_ram_n25786,
         p_wishbone_bd_ram_n25787, p_wishbone_bd_ram_n25788,
         p_wishbone_bd_ram_n25789, p_wishbone_bd_ram_n25790,
         p_wishbone_bd_ram_n25791, p_wishbone_bd_ram_n25792,
         p_wishbone_bd_ram_n25793, p_wishbone_bd_ram_n25794,
         p_wishbone_bd_ram_n25795, p_wishbone_bd_ram_n25796,
         p_wishbone_bd_ram_n25797, p_wishbone_bd_ram_n25798,
         p_wishbone_bd_ram_n25799, p_wishbone_bd_ram_n25800,
         p_wishbone_bd_ram_n25801, p_wishbone_bd_ram_n25802,
         p_wishbone_bd_ram_n25803, p_wishbone_bd_ram_n25804,
         p_wishbone_bd_ram_n25805, p_wishbone_bd_ram_n25806,
         p_wishbone_bd_ram_n25807, p_wishbone_bd_ram_n25808,
         p_wishbone_bd_ram_n25809, p_wishbone_bd_ram_n25810,
         p_wishbone_bd_ram_n25811, p_wishbone_bd_ram_n25812,
         p_wishbone_bd_ram_n25813, p_wishbone_bd_ram_n25814,
         p_wishbone_bd_ram_n25815, p_wishbone_bd_ram_n25816,
         p_wishbone_bd_ram_n25817, p_wishbone_bd_ram_n25818,
         p_wishbone_bd_ram_n25819, p_wishbone_bd_ram_n25820,
         p_wishbone_bd_ram_n25821, p_wishbone_bd_ram_n25822,
         p_wishbone_bd_ram_n25823, p_wishbone_bd_ram_n25824,
         p_wishbone_bd_ram_n25825, p_wishbone_bd_ram_n25826,
         p_wishbone_bd_ram_n25827, p_wishbone_bd_ram_n25828,
         p_wishbone_bd_ram_n25829, p_wishbone_bd_ram_n25830,
         p_wishbone_bd_ram_n25831, p_wishbone_bd_ram_n25832,
         p_wishbone_bd_ram_n25833, p_wishbone_bd_ram_n25834,
         p_wishbone_bd_ram_n25835, p_wishbone_bd_ram_n25836,
         p_wishbone_bd_ram_n25837, p_wishbone_bd_ram_n25838,
         p_wishbone_bd_ram_n25839, p_wishbone_bd_ram_n25840,
         p_wishbone_bd_ram_n25841, p_wishbone_bd_ram_n25842,
         p_wishbone_bd_ram_n25843, p_wishbone_bd_ram_n25844,
         p_wishbone_bd_ram_n25845, p_wishbone_bd_ram_n25846,
         p_wishbone_bd_ram_n25847, p_wishbone_bd_ram_n25848,
         p_wishbone_bd_ram_n25849, p_wishbone_bd_ram_n25850,
         p_wishbone_bd_ram_n25851, p_wishbone_bd_ram_n25852,
         p_wishbone_bd_ram_n25853, p_wishbone_bd_ram_n25854,
         p_wishbone_bd_ram_n25855, p_wishbone_bd_ram_n25856,
         p_wishbone_bd_ram_n25857, p_wishbone_bd_ram_n25858,
         p_wishbone_bd_ram_n25859, p_wishbone_bd_ram_n25860,
         p_wishbone_bd_ram_n25861, p_wishbone_bd_ram_n25862,
         p_wishbone_bd_ram_n25863, p_wishbone_bd_ram_n25864,
         p_wishbone_bd_ram_n25865, p_wishbone_bd_ram_n25866,
         p_wishbone_bd_ram_n25867, p_wishbone_bd_ram_n25868,
         p_wishbone_bd_ram_n25869, p_wishbone_bd_ram_n25870,
         p_wishbone_bd_ram_n25871, p_wishbone_bd_ram_n25872,
         p_wishbone_bd_ram_n25873, p_wishbone_bd_ram_n25874,
         p_wishbone_bd_ram_n25875, p_wishbone_bd_ram_n25876,
         p_wishbone_bd_ram_n25877, p_wishbone_bd_ram_n25878,
         p_wishbone_bd_ram_n25879, p_wishbone_bd_ram_n25880,
         p_wishbone_bd_ram_n25881, p_wishbone_bd_ram_n25882,
         p_wishbone_bd_ram_n25883, p_wishbone_bd_ram_n25884,
         p_wishbone_bd_ram_n25885, p_wishbone_bd_ram_n25886,
         p_wishbone_bd_ram_n25887, p_wishbone_bd_ram_n25888,
         p_wishbone_bd_ram_n25889, p_wishbone_bd_ram_n25890,
         p_wishbone_bd_ram_n25891, p_wishbone_bd_ram_n25892,
         p_wishbone_bd_ram_n25893, p_wishbone_bd_ram_n25894,
         p_wishbone_bd_ram_n25895, p_wishbone_bd_ram_n25896,
         p_wishbone_bd_ram_n25897, p_wishbone_bd_ram_n25898,
         p_wishbone_bd_ram_n25899, p_wishbone_bd_ram_n25900,
         p_wishbone_bd_ram_n25901, p_wishbone_bd_ram_n25902,
         p_wishbone_bd_ram_n25903, p_wishbone_bd_ram_n25904,
         p_wishbone_bd_ram_n25905, p_wishbone_bd_ram_n25906,
         p_wishbone_bd_ram_n25907, p_wishbone_bd_ram_n25908,
         p_wishbone_bd_ram_n25909, p_wishbone_bd_ram_n25910,
         p_wishbone_bd_ram_n25911, p_wishbone_bd_ram_n25912,
         p_wishbone_bd_ram_n25913, p_wishbone_bd_ram_n25914,
         p_wishbone_bd_ram_n25915, p_wishbone_bd_ram_n25916,
         p_wishbone_bd_ram_n25917, p_wishbone_bd_ram_n25918,
         p_wishbone_bd_ram_n25919, p_wishbone_bd_ram_n25920,
         p_wishbone_bd_ram_n25921, p_wishbone_bd_ram_n25922,
         p_wishbone_bd_ram_n25923, p_wishbone_bd_ram_n25924,
         p_wishbone_bd_ram_n25925, p_wishbone_bd_ram_n25926,
         p_wishbone_bd_ram_n25927, p_wishbone_bd_ram_n25928,
         p_wishbone_bd_ram_n25929, p_wishbone_bd_ram_n25930,
         p_wishbone_bd_ram_n25931, p_wishbone_bd_ram_n25932,
         p_wishbone_bd_ram_n25933, p_wishbone_bd_ram_n25934,
         p_wishbone_bd_ram_n25935, p_wishbone_bd_ram_n25936,
         p_wishbone_bd_ram_n25937, p_wishbone_bd_ram_n25938,
         p_wishbone_bd_ram_n25939, p_wishbone_bd_ram_n25940,
         p_wishbone_bd_ram_n25941, p_wishbone_bd_ram_n25942,
         p_wishbone_bd_ram_n25943, p_wishbone_bd_ram_n25944,
         p_wishbone_bd_ram_n25945, p_wishbone_bd_ram_n25946,
         p_wishbone_bd_ram_n25947, p_wishbone_bd_ram_n25948,
         p_wishbone_bd_ram_n25949, p_wishbone_bd_ram_n25950,
         p_wishbone_bd_ram_n25951, p_wishbone_bd_ram_n25952,
         p_wishbone_bd_ram_n25953, p_wishbone_bd_ram_n25954,
         p_wishbone_bd_ram_n25955, p_wishbone_bd_ram_n25956,
         p_wishbone_bd_ram_n25957, p_wishbone_bd_ram_n25958,
         p_wishbone_bd_ram_n25959, p_wishbone_bd_ram_n25960,
         p_wishbone_bd_ram_n25961, p_wishbone_bd_ram_n25962,
         p_wishbone_bd_ram_n25963, p_wishbone_bd_ram_n25964,
         p_wishbone_bd_ram_n25965, p_wishbone_bd_ram_n25966,
         p_wishbone_bd_ram_n25967, p_wishbone_bd_ram_n25968,
         p_wishbone_bd_ram_n25969, p_wishbone_bd_ram_n25970,
         p_wishbone_bd_ram_n25971, p_wishbone_bd_ram_n25972,
         p_wishbone_bd_ram_n25973, p_wishbone_bd_ram_n25974,
         p_wishbone_bd_ram_n25975, p_wishbone_bd_ram_n25976,
         p_wishbone_bd_ram_n25977, p_wishbone_bd_ram_n25978,
         p_wishbone_bd_ram_n25979, p_wishbone_bd_ram_n25980,
         p_wishbone_bd_ram_n25981, p_wishbone_bd_ram_n25982,
         p_wishbone_bd_ram_n25983, p_wishbone_bd_ram_n25984,
         p_wishbone_tx_fifo_N623, p_wishbone_tx_fifo_N624,
         p_wishbone_tx_fifo_N625, p_wishbone_tx_fifo_N626,
         p_wishbone_tx_fifo_N627, p_wishbone_tx_fifo_N628,
         p_wishbone_tx_fifo_N629, p_wishbone_tx_fifo_N630,
         p_wishbone_tx_fifo_N631, p_wishbone_tx_fifo_N632,
         p_wishbone_tx_fifo_N633, p_wishbone_tx_fifo_N634,
         p_wishbone_tx_fifo_N635, p_wishbone_tx_fifo_N636,
         p_wishbone_tx_fifo_N637, p_wishbone_tx_fifo_N638,
         p_wishbone_tx_fifo_N639, p_wishbone_tx_fifo_N640,
         p_wishbone_tx_fifo_N641, p_wishbone_tx_fifo_N642,
         p_wishbone_tx_fifo_N643, p_wishbone_tx_fifo_N644,
         p_wishbone_tx_fifo_N645, p_wishbone_tx_fifo_N646,
         p_wishbone_tx_fifo_N647, p_wishbone_tx_fifo_N648,
         p_wishbone_tx_fifo_N649, p_wishbone_tx_fifo_N650,
         p_wishbone_tx_fifo_N651, p_wishbone_tx_fifo_N652,
         p_wishbone_tx_fifo_N653, p_wishbone_tx_fifo_N654,
         p_wishbone_tx_fifo_n1229, p_wishbone_tx_fifo_n1230,
         p_wishbone_tx_fifo_n1231, p_wishbone_tx_fifo_n1232,
         p_wishbone_tx_fifo_n1233, p_wishbone_tx_fifo_n1234,
         p_wishbone_tx_fifo_n1235, p_wishbone_tx_fifo_n1236,
         p_wishbone_tx_fifo_n1237, p_wishbone_tx_fifo_n1238,
         p_wishbone_tx_fifo_n1239, p_wishbone_tx_fifo_n1240,
         p_wishbone_tx_fifo_n1241, p_wishbone_tx_fifo_n1242,
         p_wishbone_tx_fifo_n1243, p_wishbone_tx_fifo_n1244,
         p_wishbone_tx_fifo_n1245, p_wishbone_tx_fifo_n1246,
         p_wishbone_tx_fifo_n1247, p_wishbone_tx_fifo_n1248,
         p_wishbone_tx_fifo_n1249, p_wishbone_tx_fifo_n1250,
         p_wishbone_tx_fifo_n1251, p_wishbone_tx_fifo_n1252,
         p_wishbone_tx_fifo_n1253, p_wishbone_tx_fifo_n1254,
         p_wishbone_tx_fifo_n1255, p_wishbone_tx_fifo_n1256,
         p_wishbone_tx_fifo_n1257, p_wishbone_tx_fifo_n1258,
         p_wishbone_tx_fifo_n1259, p_wishbone_tx_fifo_n1260,
         p_wishbone_tx_fifo_n1261, p_wishbone_tx_fifo_n1262,
         p_wishbone_tx_fifo_n1263, p_wishbone_tx_fifo_n1264,
         p_wishbone_tx_fifo_n1265, p_wishbone_tx_fifo_n1266,
         p_wishbone_tx_fifo_n1267, p_wishbone_tx_fifo_n1268,
         p_wishbone_tx_fifo_n1269, p_wishbone_tx_fifo_n1270,
         p_wishbone_tx_fifo_n1271, p_wishbone_tx_fifo_n1272,
         p_wishbone_tx_fifo_n1273, p_wishbone_tx_fifo_n1274,
         p_wishbone_tx_fifo_n1275, p_wishbone_tx_fifo_n1276,
         p_wishbone_tx_fifo_n1277, p_wishbone_tx_fifo_n1278,
         p_wishbone_tx_fifo_n1279, p_wishbone_tx_fifo_n1280,
         p_wishbone_tx_fifo_n1281, p_wishbone_tx_fifo_n1282,
         p_wishbone_tx_fifo_n1283, p_wishbone_tx_fifo_n1284,
         p_wishbone_tx_fifo_n1285, p_wishbone_tx_fifo_n1286,
         p_wishbone_tx_fifo_n1287, p_wishbone_tx_fifo_n1288,
         p_wishbone_tx_fifo_n1289, p_wishbone_tx_fifo_n1290,
         p_wishbone_tx_fifo_n1291, p_wishbone_tx_fifo_n1292,
         p_wishbone_tx_fifo_n1293, p_wishbone_tx_fifo_n1294,
         p_wishbone_tx_fifo_n1295, p_wishbone_tx_fifo_n1296,
         p_wishbone_tx_fifo_n1297, p_wishbone_tx_fifo_n1298,
         p_wishbone_tx_fifo_n1299, p_wishbone_tx_fifo_n1300,
         p_wishbone_tx_fifo_n1301, p_wishbone_tx_fifo_n1302,
         p_wishbone_tx_fifo_n1303, p_wishbone_tx_fifo_n1304,
         p_wishbone_tx_fifo_n1305, p_wishbone_tx_fifo_n1306,
         p_wishbone_tx_fifo_n1307, p_wishbone_tx_fifo_n1308,
         p_wishbone_tx_fifo_n1309, p_wishbone_tx_fifo_n1310,
         p_wishbone_tx_fifo_n1311, p_wishbone_tx_fifo_n1312,
         p_wishbone_tx_fifo_n1313, p_wishbone_tx_fifo_n1314,
         p_wishbone_tx_fifo_n1315, p_wishbone_tx_fifo_n1316,
         p_wishbone_tx_fifo_n1317, p_wishbone_tx_fifo_n1318,
         p_wishbone_tx_fifo_n1319, p_wishbone_tx_fifo_n1320,
         p_wishbone_tx_fifo_n1321, p_wishbone_tx_fifo_n1322,
         p_wishbone_tx_fifo_n1323, p_wishbone_tx_fifo_n1324,
         p_wishbone_tx_fifo_n1325, p_wishbone_tx_fifo_n1326,
         p_wishbone_tx_fifo_n1327, p_wishbone_tx_fifo_n1328,
         p_wishbone_tx_fifo_n1329, p_wishbone_tx_fifo_n1330,
         p_wishbone_tx_fifo_n1331, p_wishbone_tx_fifo_n1332,
         p_wishbone_tx_fifo_n1333, p_wishbone_tx_fifo_n1334,
         p_wishbone_tx_fifo_n1335, p_wishbone_tx_fifo_n1336,
         p_wishbone_tx_fifo_n1337, p_wishbone_tx_fifo_n1338,
         p_wishbone_tx_fifo_n1339, p_wishbone_tx_fifo_n1340,
         p_wishbone_tx_fifo_n1341, p_wishbone_tx_fifo_n1342,
         p_wishbone_tx_fifo_n1343, p_wishbone_tx_fifo_n1344,
         p_wishbone_tx_fifo_n1345, p_wishbone_tx_fifo_n1346,
         p_wishbone_tx_fifo_n1347, p_wishbone_tx_fifo_n1348,
         p_wishbone_tx_fifo_n1349, p_wishbone_tx_fifo_n1350,
         p_wishbone_tx_fifo_n1351, p_wishbone_tx_fifo_n1352,
         p_wishbone_tx_fifo_n1353, p_wishbone_tx_fifo_n1354,
         p_wishbone_tx_fifo_n1355, p_wishbone_tx_fifo_n1356,
         p_wishbone_tx_fifo_n1357, p_wishbone_tx_fifo_n1358,
         p_wishbone_tx_fifo_n1359, p_wishbone_tx_fifo_n1360,
         p_wishbone_tx_fifo_n1361, p_wishbone_tx_fifo_n1362,
         p_wishbone_tx_fifo_n1363, p_wishbone_tx_fifo_n1364,
         p_wishbone_tx_fifo_n1365, p_wishbone_tx_fifo_n1366,
         p_wishbone_tx_fifo_n1367, p_wishbone_tx_fifo_n1368,
         p_wishbone_tx_fifo_n1369, p_wishbone_tx_fifo_n1370,
         p_wishbone_tx_fifo_n1371, p_wishbone_tx_fifo_n1372,
         p_wishbone_tx_fifo_n1373, p_wishbone_tx_fifo_n1374,
         p_wishbone_tx_fifo_n1375, p_wishbone_tx_fifo_n1376,
         p_wishbone_tx_fifo_n1377, p_wishbone_tx_fifo_n1378,
         p_wishbone_tx_fifo_n1379, p_wishbone_tx_fifo_n1380,
         p_wishbone_tx_fifo_n1381, p_wishbone_tx_fifo_n1382,
         p_wishbone_tx_fifo_n1383, p_wishbone_tx_fifo_n1384,
         p_wishbone_tx_fifo_n1385, p_wishbone_tx_fifo_n1386,
         p_wishbone_tx_fifo_n1387, p_wishbone_tx_fifo_n1388,
         p_wishbone_tx_fifo_n1389, p_wishbone_tx_fifo_n1390,
         p_wishbone_tx_fifo_n1391, p_wishbone_tx_fifo_n1392,
         p_wishbone_tx_fifo_n1393, p_wishbone_tx_fifo_n1394,
         p_wishbone_tx_fifo_n1395, p_wishbone_tx_fifo_n1396,
         p_wishbone_tx_fifo_n1397, p_wishbone_tx_fifo_n1398,
         p_wishbone_tx_fifo_n1399, p_wishbone_tx_fifo_n1400,
         p_wishbone_tx_fifo_n1401, p_wishbone_tx_fifo_n1402,
         p_wishbone_tx_fifo_n1403, p_wishbone_tx_fifo_n1404,
         p_wishbone_tx_fifo_n1405, p_wishbone_tx_fifo_n1406,
         p_wishbone_tx_fifo_n1407, p_wishbone_tx_fifo_n1408,
         p_wishbone_tx_fifo_n1409, p_wishbone_tx_fifo_n1410,
         p_wishbone_tx_fifo_n1411, p_wishbone_tx_fifo_n1412,
         p_wishbone_tx_fifo_n1413, p_wishbone_tx_fifo_n1414,
         p_wishbone_tx_fifo_n1415, p_wishbone_tx_fifo_n1416,
         p_wishbone_tx_fifo_n1417, p_wishbone_tx_fifo_n1418,
         p_wishbone_tx_fifo_n1419, p_wishbone_tx_fifo_n1420,
         p_wishbone_tx_fifo_n1421, p_wishbone_tx_fifo_n1422,
         p_wishbone_tx_fifo_n1423, p_wishbone_tx_fifo_n1424,
         p_wishbone_tx_fifo_n1425, p_wishbone_tx_fifo_n1426,
         p_wishbone_tx_fifo_n1427, p_wishbone_tx_fifo_n1428,
         p_wishbone_tx_fifo_n1429, p_wishbone_tx_fifo_n1430,
         p_wishbone_tx_fifo_n1431, p_wishbone_tx_fifo_n1432,
         p_wishbone_tx_fifo_n1433, p_wishbone_tx_fifo_n1434,
         p_wishbone_tx_fifo_n1435, p_wishbone_tx_fifo_n1436,
         p_wishbone_tx_fifo_n1437, p_wishbone_tx_fifo_n1438,
         p_wishbone_tx_fifo_n1439, p_wishbone_tx_fifo_n1440,
         p_wishbone_tx_fifo_n1441, p_wishbone_tx_fifo_n1442,
         p_wishbone_tx_fifo_n1443, p_wishbone_tx_fifo_n1444,
         p_wishbone_tx_fifo_n1445, p_wishbone_tx_fifo_n1446,
         p_wishbone_tx_fifo_n1447, p_wishbone_tx_fifo_n1448,
         p_wishbone_tx_fifo_n1449, p_wishbone_tx_fifo_n1450,
         p_wishbone_tx_fifo_n1451, p_wishbone_tx_fifo_n1452,
         p_wishbone_tx_fifo_n1453, p_wishbone_tx_fifo_n1454,
         p_wishbone_tx_fifo_n1455, p_wishbone_tx_fifo_n1456,
         p_wishbone_tx_fifo_n1457, p_wishbone_tx_fifo_n1458,
         p_wishbone_tx_fifo_n1459, p_wishbone_tx_fifo_n1460,
         p_wishbone_tx_fifo_n1461, p_wishbone_tx_fifo_n1462,
         p_wishbone_tx_fifo_n1463, p_wishbone_tx_fifo_n1464,
         p_wishbone_tx_fifo_n1465, p_wishbone_tx_fifo_n1466,
         p_wishbone_tx_fifo_n1467, p_wishbone_tx_fifo_n1468,
         p_wishbone_tx_fifo_n1469, p_wishbone_tx_fifo_n1470,
         p_wishbone_tx_fifo_n1471, p_wishbone_tx_fifo_n1472,
         p_wishbone_tx_fifo_n1473, p_wishbone_tx_fifo_n1474,
         p_wishbone_tx_fifo_n1475, p_wishbone_tx_fifo_n1476,
         p_wishbone_tx_fifo_n1477, p_wishbone_tx_fifo_n1478,
         p_wishbone_tx_fifo_n1479, p_wishbone_tx_fifo_n1480,
         p_wishbone_tx_fifo_n1481, p_wishbone_tx_fifo_n1482,
         p_wishbone_tx_fifo_n1483, p_wishbone_tx_fifo_n1484,
         p_wishbone_tx_fifo_n1485, p_wishbone_tx_fifo_n1486,
         p_wishbone_tx_fifo_n1487, p_wishbone_tx_fifo_n1488,
         p_wishbone_tx_fifo_n1489, p_wishbone_tx_fifo_n1490,
         p_wishbone_tx_fifo_n1491, p_wishbone_tx_fifo_n1492,
         p_wishbone_tx_fifo_n1493, p_wishbone_tx_fifo_n1494,
         p_wishbone_tx_fifo_n1495, p_wishbone_tx_fifo_n1496,
         p_wishbone_tx_fifo_n1497, p_wishbone_tx_fifo_n1498,
         p_wishbone_tx_fifo_n1499, p_wishbone_tx_fifo_n1500,
         p_wishbone_tx_fifo_n1501, p_wishbone_tx_fifo_n1502,
         p_wishbone_tx_fifo_n1503, p_wishbone_tx_fifo_n1504,
         p_wishbone_tx_fifo_n1505, p_wishbone_tx_fifo_n1506,
         p_wishbone_tx_fifo_n1507, p_wishbone_tx_fifo_n1508,
         p_wishbone_tx_fifo_n1509, p_wishbone_tx_fifo_n1510,
         p_wishbone_tx_fifo_n1511, p_wishbone_tx_fifo_n1512,
         p_wishbone_tx_fifo_n1513, p_wishbone_tx_fifo_n1514,
         p_wishbone_tx_fifo_n1515, p_wishbone_tx_fifo_n1516,
         p_wishbone_tx_fifo_n1517, p_wishbone_tx_fifo_n1518,
         p_wishbone_tx_fifo_n1519, p_wishbone_tx_fifo_n1520,
         p_wishbone_tx_fifo_n1521, p_wishbone_tx_fifo_n1522,
         p_wishbone_tx_fifo_n1523, p_wishbone_tx_fifo_n1524,
         p_wishbone_tx_fifo_n1525, p_wishbone_tx_fifo_n1526,
         p_wishbone_tx_fifo_n1527, p_wishbone_tx_fifo_n1528,
         p_wishbone_tx_fifo_n1529, p_wishbone_tx_fifo_n1530,
         p_wishbone_tx_fifo_n1531, p_wishbone_tx_fifo_n1532,
         p_wishbone_tx_fifo_n1533, p_wishbone_tx_fifo_n1534,
         p_wishbone_tx_fifo_n1535, p_wishbone_tx_fifo_n1536,
         p_wishbone_tx_fifo_n1537, p_wishbone_tx_fifo_n1538,
         p_wishbone_tx_fifo_n1539, p_wishbone_tx_fifo_n1540,
         p_wishbone_tx_fifo_n1541, p_wishbone_tx_fifo_n1542,
         p_wishbone_tx_fifo_n1543, p_wishbone_tx_fifo_n1544,
         p_wishbone_tx_fifo_n1545, p_wishbone_tx_fifo_n1546,
         p_wishbone_tx_fifo_n1547, p_wishbone_tx_fifo_n1548,
         p_wishbone_tx_fifo_n1549, p_wishbone_tx_fifo_n1550,
         p_wishbone_tx_fifo_n1551, p_wishbone_tx_fifo_n1552,
         p_wishbone_tx_fifo_n1553, p_wishbone_tx_fifo_n1554,
         p_wishbone_tx_fifo_n1555, p_wishbone_tx_fifo_n1556,
         p_wishbone_tx_fifo_n1557, p_wishbone_tx_fifo_n1558,
         p_wishbone_tx_fifo_n1559, p_wishbone_tx_fifo_n1560,
         p_wishbone_tx_fifo_n1561, p_wishbone_tx_fifo_n1562,
         p_wishbone_tx_fifo_n1563, p_wishbone_tx_fifo_n1564,
         p_wishbone_tx_fifo_n1565, p_wishbone_tx_fifo_n1566,
         p_wishbone_tx_fifo_n1567, p_wishbone_tx_fifo_n1568,
         p_wishbone_tx_fifo_n1569, p_wishbone_tx_fifo_n1570,
         p_wishbone_tx_fifo_n1571, p_wishbone_tx_fifo_n1572,
         p_wishbone_tx_fifo_n1573, p_wishbone_tx_fifo_n1574,
         p_wishbone_tx_fifo_n1575, p_wishbone_tx_fifo_n1576,
         p_wishbone_tx_fifo_n1577, p_wishbone_tx_fifo_n1578,
         p_wishbone_tx_fifo_n1579, p_wishbone_tx_fifo_n1580,
         p_wishbone_tx_fifo_n1581, p_wishbone_tx_fifo_n1582,
         p_wishbone_tx_fifo_n1583, p_wishbone_tx_fifo_n1584,
         p_wishbone_tx_fifo_n1585, p_wishbone_tx_fifo_n1586,
         p_wishbone_tx_fifo_n1587, p_wishbone_tx_fifo_n1588,
         p_wishbone_tx_fifo_n1589, p_wishbone_tx_fifo_n1590,
         p_wishbone_tx_fifo_n1591, p_wishbone_tx_fifo_n1592,
         p_wishbone_tx_fifo_n1593, p_wishbone_tx_fifo_n1594,
         p_wishbone_tx_fifo_n1595, p_wishbone_tx_fifo_n1596,
         p_wishbone_tx_fifo_n1597, p_wishbone_tx_fifo_n1598,
         p_wishbone_tx_fifo_n1599, p_wishbone_tx_fifo_n1600,
         p_wishbone_tx_fifo_n1601, p_wishbone_tx_fifo_n1602,
         p_wishbone_tx_fifo_n1603, p_wishbone_tx_fifo_n1604,
         p_wishbone_tx_fifo_n1605, p_wishbone_tx_fifo_n1606,
         p_wishbone_tx_fifo_n1607, p_wishbone_tx_fifo_n1608,
         p_wishbone_tx_fifo_n1609, p_wishbone_tx_fifo_n1610,
         p_wishbone_tx_fifo_n1611, p_wishbone_tx_fifo_n1612,
         p_wishbone_tx_fifo_n1613, p_wishbone_tx_fifo_n1614,
         p_wishbone_tx_fifo_n1615, p_wishbone_tx_fifo_n1616,
         p_wishbone_tx_fifo_n1617, p_wishbone_tx_fifo_n1618,
         p_wishbone_tx_fifo_n1619, p_wishbone_tx_fifo_n1620,
         p_wishbone_tx_fifo_n1621, p_wishbone_tx_fifo_n1622,
         p_wishbone_tx_fifo_n1623, p_wishbone_tx_fifo_n1624,
         p_wishbone_tx_fifo_n1625, p_wishbone_tx_fifo_n1626,
         p_wishbone_tx_fifo_n1627, p_wishbone_tx_fifo_n1628,
         p_wishbone_tx_fifo_n1629, p_wishbone_tx_fifo_n1630,
         p_wishbone_tx_fifo_n1631, p_wishbone_tx_fifo_n1632,
         p_wishbone_tx_fifo_n1633, p_wishbone_tx_fifo_n1634,
         p_wishbone_tx_fifo_n1635, p_wishbone_tx_fifo_n1636,
         p_wishbone_tx_fifo_n1637, p_wishbone_tx_fifo_n1638,
         p_wishbone_tx_fifo_n1639, p_wishbone_tx_fifo_n1640,
         p_wishbone_tx_fifo_n1641, p_wishbone_tx_fifo_n1642,
         p_wishbone_tx_fifo_n1643, p_wishbone_tx_fifo_n1644,
         p_wishbone_tx_fifo_n1645, p_wishbone_tx_fifo_n1646,
         p_wishbone_tx_fifo_n1647, p_wishbone_tx_fifo_n1648,
         p_wishbone_tx_fifo_n1649, p_wishbone_tx_fifo_n1650,
         p_wishbone_tx_fifo_n1651, p_wishbone_tx_fifo_n1652,
         p_wishbone_tx_fifo_n1653, p_wishbone_tx_fifo_n1654,
         p_wishbone_tx_fifo_n1655, p_wishbone_tx_fifo_n1656,
         p_wishbone_tx_fifo_n1657, p_wishbone_tx_fifo_n1658,
         p_wishbone_tx_fifo_n1659, p_wishbone_tx_fifo_n1660,
         p_wishbone_tx_fifo_n1661, p_wishbone_tx_fifo_n1662,
         p_wishbone_tx_fifo_n1663, p_wishbone_tx_fifo_n1664,
         p_wishbone_tx_fifo_n1665, p_wishbone_tx_fifo_n1666,
         p_wishbone_tx_fifo_n1667, p_wishbone_tx_fifo_n1668,
         p_wishbone_tx_fifo_n1669, p_wishbone_tx_fifo_n1670,
         p_wishbone_tx_fifo_n1671, p_wishbone_tx_fifo_n1672,
         p_wishbone_tx_fifo_n1673, p_wishbone_tx_fifo_n1674,
         p_wishbone_tx_fifo_n1675, p_wishbone_tx_fifo_n1676,
         p_wishbone_tx_fifo_n1677, p_wishbone_tx_fifo_n1678,
         p_wishbone_tx_fifo_n1679, p_wishbone_tx_fifo_n1680,
         p_wishbone_tx_fifo_n1681, p_wishbone_tx_fifo_n1682,
         p_wishbone_tx_fifo_n1683, p_wishbone_tx_fifo_n1684,
         p_wishbone_tx_fifo_n1685, p_wishbone_tx_fifo_n1686,
         p_wishbone_tx_fifo_n1687, p_wishbone_tx_fifo_n1688,
         p_wishbone_tx_fifo_n1689, p_wishbone_tx_fifo_n1690,
         p_wishbone_tx_fifo_n1691, p_wishbone_tx_fifo_n1692,
         p_wishbone_tx_fifo_n1693, p_wishbone_tx_fifo_n1694,
         p_wishbone_tx_fifo_n1695, p_wishbone_tx_fifo_n1696,
         p_wishbone_tx_fifo_n1697, p_wishbone_tx_fifo_n1698,
         p_wishbone_tx_fifo_n1699, p_wishbone_tx_fifo_n1700,
         p_wishbone_tx_fifo_n1701, p_wishbone_tx_fifo_n1702,
         p_wishbone_tx_fifo_n1703, p_wishbone_tx_fifo_n1704,
         p_wishbone_tx_fifo_n1705, p_wishbone_tx_fifo_n1706,
         p_wishbone_tx_fifo_n1707, p_wishbone_tx_fifo_n1708,
         p_wishbone_tx_fifo_n1709, p_wishbone_tx_fifo_n1710,
         p_wishbone_tx_fifo_n1711, p_wishbone_tx_fifo_n1712,
         p_wishbone_tx_fifo_n1713, p_wishbone_tx_fifo_n1714,
         p_wishbone_tx_fifo_n1715, p_wishbone_tx_fifo_n1716,
         p_wishbone_tx_fifo_n1717, p_wishbone_tx_fifo_n1718,
         p_wishbone_tx_fifo_n1719, p_wishbone_tx_fifo_n1720,
         p_wishbone_tx_fifo_n1721, p_wishbone_tx_fifo_n1722,
         p_wishbone_tx_fifo_n1723, p_wishbone_tx_fifo_n1724,
         p_wishbone_tx_fifo_n1725, p_wishbone_tx_fifo_n1726,
         p_wishbone_tx_fifo_n1727, p_wishbone_tx_fifo_n1728,
         p_wishbone_tx_fifo_n1729, p_wishbone_tx_fifo_n1730,
         p_wishbone_tx_fifo_n1731, p_wishbone_tx_fifo_n1732,
         p_wishbone_tx_fifo_n1733, p_wishbone_tx_fifo_n1734,
         p_wishbone_tx_fifo_n1735, p_wishbone_tx_fifo_n1736,
         p_wishbone_tx_fifo_n1737, p_wishbone_tx_fifo_n1738,
         p_wishbone_tx_fifo_n1739, p_wishbone_tx_fifo_n1740,
         p_wishbone_tx_fifo_n1741, p_wishbone_tx_fifo_n1742,
         p_wishbone_tx_fifo_n1743, p_wishbone_tx_fifo_n1744,
         p_wishbone_tx_fifo_n1745, p_wishbone_tx_fifo_n1746,
         p_wishbone_tx_fifo_n1747, p_wishbone_tx_fifo_n1748,
         p_wishbone_tx_fifo_n1749, p_wishbone_tx_fifo_n1750,
         p_wishbone_tx_fifo_n1751, p_wishbone_tx_fifo_n1752,
         p_wishbone_tx_fifo_n1753, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35897, n33925, n35892, n33930, n35893,
         n35894, n33926, n35895, n35896, n35885, n35886, n35887, n35888,
         n35889, n35890, n35884, n35891, n35883, n35882, n35877, n35878,
         n35879, n35880, n35881, p_rxethmac1_crcrx_N25, p_rxethmac1_crcrx_N21,
         p_rxethmac1_crcrx_N17, p_rxethmac1_crcrx_N13, p_rxethmac1_crcrx_N9,
         p_rxethmac1_crcrx_N5, p_rxethmac1_crcrx_N8, p_rxethmac1_crcrx_N26,
         p_rxethmac1_crcrx_N22, p_rxethmac1_crcrx_N18, p_rxethmac1_crcrx_N14,
         p_rxethmac1_crcrx_N10, p_rxethmac1_crcrx_N6, p_rxethmac1_crcrx_N34,
         p_rxethmac1_crcrx_N30, p_rxethmac1_crcrx_N4, p_rxethmac1_crcrx_N32,
         p_rxethmac1_crcrx_N28, p_rxethmac1_crcrx_N24, p_rxethmac1_crcrx_N20,
         p_rxethmac1_crcrx_N16, p_rxethmac1_crcrx_N12, p_rxethmac1_crcrx_N33,
         p_rxethmac1_crcrx_N29, p_rxethmac1_crcrx_N31, p_rxethmac1_crcrx_N27,
         p_rxethmac1_crcrx_N23, p_rxethmac1_crcrx_N19, p_rxethmac1_crcrx_N15,
         p_rxethmac1_crcrx_N11, p_rxethmac1_crcrx_N7, p_rxethmac1_crcrx_N3,
         p_wishbone_rx_fifo_N623, p_wishbone_rx_fifo_N624,
         p_wishbone_rx_fifo_N625, p_wishbone_rx_fifo_N626,
         p_wishbone_rx_fifo_N627, p_wishbone_rx_fifo_N628,
         p_wishbone_rx_fifo_N629, p_wishbone_rx_fifo_N630,
         p_wishbone_rx_fifo_N631, p_wishbone_rx_fifo_N632,
         p_wishbone_rx_fifo_N633, p_wishbone_rx_fifo_N634,
         p_wishbone_rx_fifo_N635, p_wishbone_rx_fifo_N636,
         p_wishbone_rx_fifo_N637, p_wishbone_rx_fifo_N638,
         p_wishbone_rx_fifo_N639, p_wishbone_rx_fifo_N640,
         p_wishbone_rx_fifo_N641, p_wishbone_rx_fifo_N642,
         p_wishbone_rx_fifo_N643, p_wishbone_rx_fifo_N644,
         p_wishbone_rx_fifo_N645, p_wishbone_rx_fifo_N646,
         p_wishbone_rx_fifo_N647, p_wishbone_rx_fifo_N648,
         p_wishbone_rx_fifo_N649, p_wishbone_rx_fifo_N650,
         p_wishbone_rx_fifo_N651, p_wishbone_rx_fifo_N652,
         p_wishbone_rx_fifo_N653, p_wishbone_rx_fifo_N654, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468;
  wire   n31339, n31354, n31365, n31377, n31388, n32001, n64123, n64122,
         n64461, n56483, n56485, n56478, n56396, n56464, n56460, n56459,
         n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404,
         n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56394,
         n56413, n56414, n56470, n56416, n56418, n56419, n56420, n56421,
         n56438, n56427, n56426, n56424, n56423, n56422, n56430, n56437,
         n56435, n56462, n56372, n56440, n56486, n56457, n56456, n56455,
         n56454, n56453, n56452, n56451, n56450, n56449, n56448, n56447,
         n56446, n56445, n56444, n56443, n56377, n56376, n56375, n56374,
         n56373, n56442, n56393, n56388, n56387, n56381, n56370, n56369,
         n56368, n56367, n56366, n56365, n56364, n56363, n56362, n56361,
         n56360, n56359, n56358, n56357, n56356, n56355, n56354, n56353,
         n56352, n56351, n56350, n56349, n56348, n56347, n56346, n56345,
         n56344, n56343, n56342, n56371, n56340, n56339, n56338, n56337,
         n56336, n56335, n56334, n56333, n56332, n56331, n56330, n56329,
         n56328, n56327, n56326, n56325, n56324, n56323, n56322, n56321,
         n56320, n56319, n56318, n56317, n56316, n56315, n56314, n56313,
         n56312, n56341, n56311, n64121, n64119, n64116, n64114, n64113,
         n64111, n64108, n64106, n64105, n64103, n64100, n64098, n64097,
         n64095, n64092, n64090, n64089, n64087, n64084, n64082, n64081,
         n64079, n64076, n64074, n64073, n64071, n64068, n64066, n64065,
         n64063, n64060, n64058, n64057, n64055, n64052, n64050, n64049,
         n64047, n64044, n64042, n64041, n64039, n64036, n64034, n64033,
         n64031, n64028, n64026, n64025, n64023, n64020, n64018, n64017,
         n64015, n64012, n64010, n64009, n64007, n64004, n64002, n64001,
         n63999, n63996, n63994, n63993, n63991, n63988, n63986, n63985,
         n63983, n63980, n63978, n63977, n63975, n63972, n63970, n63969,
         n63967, n63964, n63962, n63961, n63959, n63956, n63954, n63953,
         n63951, n63948, n63946, n63945, n63943, n63940, n63938, n63937,
         n63935, n63932, n63930, n63929, n63927, n63924, n63922, n63921,
         n63919, n63916, n63914, n63913, n63911, n63908, n63906, n63905,
         n63903, n63900, n63898, n63897, n63895, n63892, n63890, n63889,
         n63887, n63884, n63882, n63881, n63879, n63876, n63874, n63873,
         n63871, n63868, n63866, n63865, n63863, n63860, n63858, n63857,
         n63855, n63852, n63850, n63849, n63847, n63844, n63842, n63841,
         n63839, n63836, n63834, n63833, n63831, n63828, n63826, n63825,
         n63823, n63820, n63818, n63817, n63815, n63812, n63810, n63809,
         n63807, n63804, n63802, n63801, n63799, n63796, n63794, n63793,
         n63791, n63788, n63786, n63785, n63783, n63780, n63778, n63777,
         n63775, n63772, n63770, n63769, n63767, n63764, n63762, n63761,
         n63759, n63756, n63754, n63753, n63751, n63748, n63746, n63745,
         n63743, n63740, n63738, n63737, n63735, n63732, n63730, n63729,
         n63727, n63724, n63722, n63721, n63719, n63716, n63714, n63713,
         n63711, n63708, n63706, n63705, n63703, n63700, n63698, n63697,
         n63695, n63692, n63690, n63689, n63687, n63684, n63682, n63681,
         n63679, n63676, n63674, n63673, n63671, n63668, n63666, n63665,
         n63663, n63660, n63658, n63657, n63655, n63652, n63650, n63649,
         n63647, n63644, n63642, n63641, n63639, n63636, n63634, n63633,
         n63631, n63628, n63626, n63625, n63623, n63620, n63618, n63617,
         n63615, n63612, n63610, n63609, n63607, n63604, n63602, n63601,
         n63599, n63596, n63594, n63593, n63591, n63588, n63586, n63585,
         n63583, n63580, n63578, n63577, n63575, n63572, n63570, n63569,
         n63567, n63564, n63562, n63561, n63559, n63556, n63554, n63553,
         n63551, n63548, n63546, n63545, n63543, n63540, n63538, n63537,
         n63535, n63532, n63530, n63529, n63527, n63524, n63522, n63521,
         n63519, n63516, n63514, n63513, n63511, n63508, n63506, n63505,
         n63503, n63500, n63498, n63497, n63496, n63495, n63494, n63493,
         n63491, n63488, n63486, n63485, n63483, n63480, n63478, n63477,
         n63475, n63472, n63470, n63469, n63467, n63464, n63462, n63461,
         n63459, n63456, n63454, n63449, n63447, n63444, n63442, n63441,
         n63439, n63436, n63434, n63433, n63431, n63428, n63426, n63425,
         n63423, n63420, n63418, n63417, n63415, n63412, n63410, n63409,
         n63408, n63407, n63406, n63405, n63403, n63400, n63398, n63397,
         n63395, n63392, n63390, n63389, n63387, n63384, n63382, n63381,
         n63379, n63376, n63374, n63373, n63371, n63368, n63366, n63365,
         n63363, n63360, n63358, n63357, n63356, n63355, n63354, n63353,
         n63351, n63348, n63346, n63345, n63343, n63340, n63338, n63337,
         n63335, n63332, n63330, n63329, n63327, n63324, n63322, n63321,
         n63319, n63316, n63314, n63313, n63311, n63308, n63306, n63305,
         n63303, n63300, n63298, n63297, n63295, n63292, n63290, n63289,
         n63288, n63287, n63286, n63285, n63283, n63280, n63278, n63277,
         n63275, n63272, n63270, n63269, n63267, n63264, n63262, n63261,
         n63259, n63256, n63254, n63253, n63251, n63248, n63246, n63245,
         n63243, n63240, n63238, n63237, n63235, n63232, n63230, n63229,
         n63227, n63224, n63222, n63221, n63219, n63216, n63214, n63213,
         n63211, n63208, n63206, n63205, n63203, n63200, n63198, n63197,
         n63195, n63192, n63190, n63189, n63187, n63184, n63182, n63181,
         n63179, n63176, n63174, n63173, n63171, n63168, n63166, n63165,
         n63163, n63160, n63158, n63157, n63156, n63155, n63154, n63153,
         n63152, n63151, n63150, n63149, n63147, n63144, n63142, n63141,
         n63139, n63136, n63134, n63133, n63132, n63131, n63130, n63129,
         n63127, n63124, n63122, n63121, n63119, n63116, n63114, n63113,
         n63111, n63108, n63106, n63105, n63103, n63100, n63098, n63097,
         n63095, n63092, n63090, n63089, n63088, n63087, n63086, n63085,
         n63083, n63080, n63078, n63077, n63075, n63072, n63070, n63069,
         n63068, n63067, n63066, n63065, n63063, n63060, n63058, n63057,
         n63055, n63052, n63050, n63049, n63047, n63044, n63042, n63041,
         n63039, n63036, n63034, n63033, n63031, n63028, n63026, n63025,
         n63023, n63020, n63018, n63017, n63015, n63012, n63010, n63009,
         n63008, n63007, n63006, n63005, n63004, n63003, n63002, n63001,
         n62999, n62996, n62994, n62993, n62992, n62991, n62990, n62989,
         n62987, n62984, n62982, n62981, n62979, n62976, n62974, n62973,
         n62971, n62968, n62966, n62965, n62963, n62960, n62958, n62957,
         n62956, n62955, n62954, n62953, n62951, n62948, n62946, n62945,
         n62943, n62940, n62938, n62937, n62935, n62932, n62930, n62929,
         n62927, n62924, n62922, n62921, n62919, n62916, n62914, n62913,
         n62911, n62908, n62906, n62905, n62903, n62900, n62898, n62897,
         n62896, n62895, n62894, n62893, n62891, n62888, n62886, n62885,
         n62883, n62880, n62878, n62877, n62876, n62875, n62874, n62873,
         n62871, n62868, n62866, n62865, n62863, n62860, n62858, n62857,
         n62855, n62852, n62850, n62849, n62847, n62844, n62842, n62841,
         n62839, n62836, n62834, n62833, n62831, n62828, n62826, n62825,
         n62823, n62820, n62818, n62817, n62815, n62812, n62810, n62809,
         n62808, n62807, n62806, n62805, n62803, n62800, n62798, n62797,
         n62795, n62792, n62790, n62789, n62788, n62787, n62786, n62785,
         n62783, n62780, n62778, n62777, n62775, n62772, n62770, n62769,
         n62767, n62764, n62762, n62761, n62759, n62756, n62754, n62753,
         n62751, n62748, n62746, n62745, n62743, n62740, n62738, n62737,
         n62736, n62735, n62734, n62733, n62732, n62731, n62730, n62729,
         n62727, n62724, n62722, n62721, n62719, n62716, n62714, n62713,
         n62711, n62708, n62706, n62705, n62703, n62700, n62698, n62697,
         n62695, n62692, n62690, n62689, n62687, n62684, n62682, n62681,
         n62679, n62676, n62674, n62673, n62671, n62668, n62666, n62665,
         n62663, n62660, n62658, n62657, n62655, n62652, n62650, n62649,
         n62647, n62644, n62642, n62641, n62639, n62636, n62634, n62633,
         n62631, n62628, n62626, n62625, n62623, n62620, n62618, n62617,
         n62615, n62612, n62610, n62609, n62607, n62604, n62602, n62601,
         n62599, n62596, n62594, n62593, n62591, n62588, n62586, n62585,
         n62584, n62583, n62582, n62581, n62579, n62576, n62574, n62569,
         n62567, n62564, n62562, n62561, n62559, n62556, n62554, n62553,
         n62551, n62548, n62546, n62545, n62543, n62540, n62538, n62537,
         n62535, n62532, n62530, n62529, n62527, n62524, n62522, n62517,
         n62515, n62512, n62510, n62509, n62507, n62504, n62502, n62501,
         n62499, n62496, n62494, n62493, n62492, n62491, n62490, n62489,
         n62487, n62484, n62482, n62481, n62479, n62476, n62474, n62473,
         n62471, n62468, n62466, n62465, n62463, n62460, n62458, n62457,
         n62455, n62452, n62450, n62449, n62447, n62444, n62442, n62441,
         n62439, n62436, n62434, n62429, n62427, n62424, n62422, n62421,
         n62420, n62419, n62418, n62417, n62416, n62415, n62414, n62413,
         n62412, n62411, n62410, n62409, n62407, n62404, n62402, n62401,
         n62399, n62396, n62394, n62393, n62391, n62388, n62386, n62385,
         n62384, n62383, n62382, n62381, n62379, n62376, n62374, n62369,
         n62367, n62364, n62362, n62357, n62355, n62352, n62350, n62349,
         n62348, n62347, n62346, n62333, n62332, n62331, n62330, n62329,
         n62327, n62324, n62322, n62321, n62319, n62316, n62314, n62313,
         n62311, n62308, n62306, n62305, n62304, n62303, n62302, n62301,
         n62299, n62296, n62294, n62293, n62291, n62288, n62286, n62285,
         n62284, n62283, n62282, n62281, n62280, n62279, n62278, n62277,
         n62275, n62272, n62270, n62269, n62267, n62264, n62262, n62261,
         n62259, n62256, n62254, n62253, n62251, n62248, n62246, n62245,
         n62243, n62240, n62238, n62237, n62235, n62232, n62230, n62229,
         n62227, n62224, n62222, n62221, n62219, n62216, n62214, n62213,
         n62211, n62208, n62206, n62205, n62203, n62200, n62198, n62197,
         n62195, n62192, n62190, n62189, n62187, n62184, n62182, n62181,
         n62179, n62176, n62174, n62173, n62171, n62168, n62166, n62165,
         n62163, n62160, n62158, n62157, n62155, n62152, n62150, n62149,
         n62147, n62144, n62142, n62141, n62139, n62136, n62134, n62133,
         n62131, n62128, n62126, n62125, n62123, n62120, n62118, n62117,
         n62115, n62112, n62110, n62109, n62107, n62104, n62102, n62101,
         n62099, n62096, n62094, n62093, n62091, n62088, n62086, n62085,
         n62083, n62080, n62078, n62077, n62075, n62072, n62070, n62069,
         n62067, n62064, n62062, n62061, n62059, n62056, n62054, n62053,
         n62051, n62048, n62046, n62045, n62043, n62040, n62038, n62037,
         n62035, n62032, n62030, n62029, n62027, n62024, n62022, n62021,
         n62019, n62016, n62014, n62013, n62011, n62008, n62006, n62005,
         n62003, n62000, n61998, n61997, n61995, n61992, n61990, n61989,
         n61987, n61984, n61982, n61981, n61979, n61976, n61974, n61973,
         n61971, n61968, n61966, n61965, n61963, n61960, n61958, n61957,
         n61955, n61952, n61950, n61949, n61947, n61944, n61942, n61941,
         n61939, n61936, n61934, n61933, n61931, n61928, n61926, n61925,
         n61923, n61920, n61918, n61917, n61915, n61912, n61910, n61909,
         n61907, n61904, n61902, n61901, n61899, n61896, n61894, n61893,
         n61891, n61888, n61886, n61885, n61883, n61880, n61878, n61877,
         n61875, n61872, n61870, n61869, n61867, n61864, n61862, n61861,
         n61859, n61856, n61854, n61853, n61851, n61848, n61846, n61845,
         n61843, n61840, n61838, n61837, n61835, n61832, n61830, n61829,
         n61827, n61824, n61822, n61821, n61819, n61816, n61814, n61813,
         n61811, n61808, n61806, n61805, n61803, n61800, n61798, n61797,
         n61795, n61792, n61790, n61789, n61787, n61784, n61782, n61781,
         n61779, n61776, n61774, n61773, n61771, n61768, n61766, n61765,
         n61763, n61760, n61758, n61757, n61755, n61752, n61750, n61749,
         n61747, n61744, n61742, n61741, n61739, n61736, n61734, n61733,
         n61731, n61728, n61726, n61725, n61723, n61720, n61718, n61717,
         n61715, n61712, n61710, n61709, n61707, n61704, n61702, n61701,
         n61699, n61696, n61694, n61693, n61691, n61688, n61686, n61685,
         n61683, n61680, n61678, n61677, n61675, n61672, n61670, n61669,
         n61667, n61664, n61662, n61661, n61659, n61656, n61654, n61653,
         n61651, n61648, n61646, n61645, n61643, n61640, n61638, n61637,
         n61635, n61632, n61630, n61629, n61627, n61624, n61622, n61621,
         n61619, n61616, n61614, n61613, n61611, n61608, n61606, n61605,
         n61604, n61603, n61602, n61601, n61599, n61596, n61594, n61593,
         n61591, n61588, n61586, n61585, n61583, n61580, n61578, n61577,
         n61575, n61572, n61570, n61569, n61567, n61564, n61562, n61557,
         n61555, n61552, n61550, n61549, n61547, n61544, n61542, n61541,
         n61539, n61536, n61534, n61533, n61531, n61528, n61526, n61525,
         n61523, n61520, n61518, n61517, n61516, n61515, n61514, n61513,
         n61511, n61508, n61506, n61505, n61503, n61500, n61498, n61497,
         n61495, n61492, n61490, n61489, n61487, n61484, n61482, n61481,
         n61479, n61476, n61474, n61473, n61471, n61468, n61466, n61465,
         n61464, n61463, n61462, n61461, n61459, n61456, n61454, n61453,
         n61451, n61448, n61446, n61445, n61443, n61440, n61438, n61437,
         n61435, n61432, n61430, n61429, n61427, n61424, n61422, n61421,
         n61419, n61416, n61414, n61413, n61411, n61408, n61406, n61405,
         n61403, n61400, n61398, n61397, n61396, n61395, n61394, n61393,
         n61391, n61388, n61386, n61385, n61383, n61380, n61378, n61377,
         n61375, n61372, n61370, n61369, n61367, n61364, n61362, n61361,
         n61359, n61356, n61354, n61353, n61351, n61348, n61346, n61345,
         n61343, n61340, n61338, n61337, n61336, n61335, n61334, n61333,
         n61331, n61328, n61326, n61325, n61323, n61320, n61318, n61317,
         n61315, n61312, n61310, n61309, n61307, n61304, n61302, n61301,
         n61299, n61296, n61294, n61293, n61292, n61291, n61290, n61289,
         n61287, n61284, n61282, n61281, n61279, n61276, n61274, n61273,
         n61272, n61271, n61270, n61269, n61267, n61264, n61262, n61261,
         n61259, n61256, n61254, n61253, n61251, n61248, n61246, n61245,
         n61243, n61240, n61238, n61237, n61235, n61232, n61230, n61229,
         n61227, n61224, n61222, n61221, n61219, n61216, n61214, n61213,
         n61212, n61211, n61210, n61209, n61208, n61207, n61206, n61205,
         n61203, n61200, n61198, n61197, n61196, n61195, n61194, n61193,
         n61191, n61188, n61186, n61185, n61183, n61180, n61178, n61177,
         n61175, n61172, n61170, n61169, n61167, n61164, n61162, n61161,
         n61160, n61159, n61158, n61157, n61155, n61152, n61150, n61149,
         n61147, n61144, n61142, n61141, n61139, n61136, n61134, n61133,
         n61131, n61128, n61126, n61125, n61123, n61120, n61118, n61117,
         n61115, n61112, n61110, n61109, n61107, n61104, n61102, n61101,
         n61100, n61099, n61098, n61097, n61095, n61092, n61090, n61089,
         n61087, n61084, n61082, n61081, n61080, n61079, n61078, n61077,
         n61075, n61072, n61070, n61069, n61067, n61064, n61062, n61061,
         n61059, n61056, n61054, n61053, n61051, n61048, n61046, n61045,
         n61043, n61040, n61038, n61037, n61035, n61032, n61030, n61029,
         n61027, n61024, n61022, n61021, n61019, n61016, n61014, n61013,
         n61012, n61011, n61010, n61009, n61007, n61004, n61002, n61001,
         n60999, n60996, n60994, n60993, n60992, n60991, n60990, n60989,
         n60987, n60984, n60982, n60981, n60979, n60976, n60974, n60973,
         n60971, n60968, n60966, n60965, n60963, n60960, n60958, n60957,
         n60955, n60952, n60950, n60949, n60947, n60944, n60942, n60941,
         n60940, n60939, n60938, n60937, n60936, n60935, n60934, n60933,
         n60931, n60928, n60926, n60925, n60923, n60920, n60918, n60917,
         n60915, n60912, n60910, n60909, n60907, n60904, n60902, n60901,
         n60899, n60896, n60894, n60893, n60891, n60888, n60886, n60885,
         n60883, n60880, n60878, n60877, n60875, n60872, n60870, n60869,
         n60867, n60864, n60862, n60861, n60859, n60856, n60854, n60853,
         n60851, n60848, n60846, n60845, n60843, n60840, n60838, n60837,
         n60835, n60832, n60830, n60829, n60827, n60824, n60822, n60821,
         n60819, n60816, n60814, n60813, n60811, n60808, n60806, n60805,
         n60804, n60803, n60802, n60801, n60800, n60799, n60798, n60797,
         n60795, n60792, n60790, n60789, n60787, n60784, n60782, n60781,
         n60779, n60776, n60774, n60773, n60771, n60768, n60766, n60765,
         n60763, n60760, n60758, n60757, n60755, n60752, n60750, n60749,
         n60747, n60744, n60742, n60741, n60739, n60736, n60734, n60733,
         n60731, n60728, n60726, n60725, n60723, n60720, n60718, n60717,
         n60715, n60712, n60710, n60709, n60707, n60704, n60702, n60701,
         n60700, n60699, n60698, n60697, n60695, n60692, n60690, n60689,
         n60688, n60687, n60686, n60685, n60683, n60680, n60678, n60677,
         n60675, n60672, n60670, n60669, n60667, n60664, n60662, n60661,
         n60659, n60656, n60654, n60653, n60651, n60648, n60646, n60645,
         n60644, n60643, n60642, n60641, n60639, n60636, n60634, n60633,
         n60631, n60628, n60626, n60625, n60623, n60620, n60618, n60617,
         n60616, n60615, n60614, n60613, n60611, n60608, n60606, n60605,
         n60603, n60600, n60598, n60597, n60596, n60595, n60594, n60593,
         n60591, n60588, n60586, n60585, n60583, n60580, n60578, n60577,
         n60575, n60572, n60570, n60569, n60567, n60564, n60562, n60561,
         n60560, n60559, n60558, n60557, n60555, n60552, n60550, n60545,
         n60544, n60543, n60542, n60541, n60540, n60539, n60538, n60537,
         n60535, n60532, n60530, n60529, n60527, n60524, n60522, n60521,
         n60520, n60519, n60518, n60517, n60516, n60515, n60514, n60513,
         n60512, n60511, n60510, n60509, n60507, n60504, n60502, n60501,
         n60500, n60499, n60498, n60497, n60495, n60492, n60490, n60489,
         n60488, n60487, n60486, n60485, n60483, n60480, n60478, n60477,
         n60476, n60475, n60474, n60473, n60472, n60471, n60470, n60469,
         n60467, n60464, n60462, n60453, n60451, n60448, n60446, n60445,
         n60443, n60440, n60438, n60437, n60435, n60432, n60430, n60429,
         n60428, n60427, n60426, n60425, n60423, n60420, n60418, n60417,
         n60415, n60412, n60410, n60409, n60407, n60404, n60402, n60401,
         n60399, n60396, n60394, n60393, n60391, n60388, n60386, n60385,
         n60383, n60380, n60378, n60377, n60375, n60372, n60370, n60369,
         n60367, n60364, n60362, n60361, n60359, n60356, n60354, n60353,
         n60351, n60348, n60346, n60345, n60343, n60340, n60338, n60337,
         n60335, n60332, n60330, n60329, n60327, n60324, n60322, n60321,
         n60319, n60316, n60314, n60313, n60311, n60308, n60306, n60305,
         n60303, n60300, n60298, n60297, n60295, n60292, n60290, n60289,
         n60287, n60284, n60282, n60281, n60279, n60276, n60274, n60273,
         n60271, n60268, n60266, n60265, n60263, n60260, n60258, n60257,
         n60255, n60252, n60250, n60249, n60247, n60244, n60242, n60241,
         n60239, n60236, n60234, n60233, n60231, n60228, n60226, n60225,
         n60223, n60220, n60218, n60217, n60215, n60212, n60210, n60209,
         n60207, n60204, n60202, n60201, n60199, n60196, n60194, n60193,
         n60191, n60188, n60186, n60185, n60183, n60180, n60178, n60177,
         n60175, n60172, n60170, n60169, n60167, n60164, n60162, n60161,
         n60159, n60156, n60154, n60153, n60151, n60148, n60146, n60145,
         n60143, n60140, n60138, n60137, n60135, n60132, n60130, n60129,
         n60127, n60124, n60122, n60121, n60119, n60116, n60114, n60113,
         n60111, n60108, n60106, n60105, n60103, n60100, n60098, n60097,
         n60095, n60092, n60090, n60089, n60087, n60084, n60082, n60081,
         n60079, n60076, n60074, n60073, n60071, n60068, n60066, n60065,
         n60063, n60060, n60058, n60057, n60055, n60052, n60050, n60049,
         n60047, n60044, n60042, n60041, n60039, n60036, n60034, n60033,
         n60031, n60028, n60026, n60025, n60023, n60020, n60018, n60017,
         n60015, n60012, n60010, n60009, n60007, n60004, n60002, n60001,
         n59999, n59996, n59994, n59993, n59991, n59988, n59986, n59985,
         n59983, n59980, n59978, n59977, n59975, n59972, n59970, n59969,
         n59967, n59964, n59962, n59961, n59959, n59956, n59954, n59953,
         n59951, n59948, n59946, n59945, n59943, n59940, n59938, n59937,
         n59935, n59932, n59930, n59929, n59927, n59924, n59922, n59921,
         n59919, n59916, n59914, n59913, n59911, n59908, n59906, n59905,
         n59903, n59900, n59898, n59897, n59895, n59892, n59890, n59889,
         n59887, n59884, n59882, n59881, n59879, n59876, n59874, n59873,
         n59871, n59868, n59866, n59865, n59863, n59860, n59858, n59857,
         n59855, n59852, n59850, n59849, n59847, n59844, n59842, n59841,
         n59839, n59836, n59834, n59833, n59831, n59828, n59826, n59825,
         n59823, n59820, n59818, n59817, n59815, n59812, n59810, n59809,
         n59807, n59804, n59802, n59801, n59799, n59796, n59794, n59793,
         n59791, n59788, n59786, n59785, n59783, n59780, n59778, n59777,
         n59775, n59772, n59770, n59769, n59767, n59764, n59762, n59761,
         n59759, n59756, n59754, n59753, n59751, n59748, n59746, n59745,
         n59743, n59740, n59738, n59737, n59735, n59732, n59730, n59729,
         n59727, n59724, n59722, n59721, n59719, n59716, n59714, n59713,
         n59712, n59711, n59710, n59709, n59707, n59704, n59702, n59701,
         n59699, n59696, n59694, n59693, n59691, n59688, n59686, n59685,
         n59683, n59680, n59678, n59677, n59675, n59672, n59670, n59665,
         n59663, n59660, n59658, n59657, n59655, n59652, n59650, n59649,
         n59647, n59644, n59642, n59641, n59639, n59636, n59634, n59633,
         n59631, n59628, n59626, n59625, n59624, n59623, n59622, n59621,
         n59619, n59616, n59614, n59613, n59611, n59608, n59606, n59605,
         n59603, n59600, n59598, n59597, n59595, n59592, n59590, n59589,
         n59587, n59584, n59582, n59581, n59579, n59576, n59574, n59573,
         n59572, n59571, n59570, n59569, n59567, n59564, n59562, n59561,
         n59559, n59556, n59554, n59553, n59551, n59548, n59546, n59545,
         n59543, n59540, n59538, n59537, n59535, n59532, n59530, n59529,
         n59527, n59524, n59522, n59521, n59519, n59516, n59514, n59513,
         n59511, n59508, n59506, n59505, n59504, n59503, n59502, n59501,
         n59499, n59496, n59494, n59493, n59491, n59488, n59486, n59485,
         n59483, n59480, n59478, n59477, n59475, n59472, n59470, n59469,
         n59467, n59464, n59462, n59461, n59459, n59456, n59454, n59453,
         n59451, n59448, n59446, n59445, n59444, n59443, n59442, n59441,
         n59439, n59436, n59434, n59433, n59431, n59428, n59426, n59425,
         n59423, n59420, n59418, n59417, n59415, n59412, n59410, n59409,
         n59407, n59404, n59402, n59401, n59400, n59399, n59398, n59397,
         n59395, n59392, n59390, n59389, n59387, n59384, n59382, n59381,
         n59380, n59379, n59378, n59377, n59375, n59372, n59370, n59369,
         n59367, n59364, n59362, n59361, n59359, n59356, n59354, n59353,
         n59351, n59348, n59346, n59345, n59343, n59340, n59338, n59337,
         n59335, n59332, n59330, n59329, n59327, n59324, n59322, n59321,
         n59320, n59319, n59318, n59317, n59316, n59315, n59314, n59313,
         n59311, n59308, n59306, n59305, n59304, n59303, n59302, n59301,
         n59299, n59296, n59294, n59293, n59291, n59288, n59286, n59285,
         n59283, n59280, n59278, n59277, n59275, n59272, n59270, n59269,
         n59268, n59267, n59266, n59265, n59263, n59260, n59258, n59257,
         n59255, n59252, n59250, n59249, n59247, n59244, n59242, n59241,
         n59239, n59236, n59234, n59233, n59231, n59228, n59226, n59225,
         n59223, n59220, n59218, n59217, n59215, n59212, n59210, n59209,
         n59208, n59207, n59206, n59205, n59203, n59200, n59198, n59197,
         n59195, n59192, n59190, n59189, n59188, n59187, n59186, n59185,
         n59183, n59180, n59178, n59177, n59175, n59172, n59170, n59169,
         n59167, n59164, n59162, n59161, n59159, n59156, n59154, n59153,
         n59151, n59148, n59146, n59145, n59143, n59140, n59138, n59137,
         n59135, n59132, n59130, n59129, n59127, n59124, n59122, n59121,
         n59120, n59119, n59118, n59117, n59115, n59112, n59110, n59109,
         n59107, n59104, n59102, n59101, n59100, n59099, n59098, n59097,
         n59095, n59092, n59090, n59089, n59087, n59084, n59082, n59081,
         n59079, n59076, n59074, n59073, n59071, n59068, n59066, n59065,
         n59063, n59060, n59058, n59057, n59055, n59052, n59050, n59049,
         n59048, n59047, n59046, n59045, n59044, n59043, n59042, n59041,
         n59039, n59036, n59034, n59033, n59031, n59028, n59026, n59025,
         n59023, n59020, n59018, n59017, n59015, n59012, n59010, n59009,
         n59007, n59004, n59002, n59001, n58999, n58996, n58994, n58993,
         n58991, n58988, n58986, n58985, n58983, n58980, n58978, n58977,
         n58975, n58972, n58970, n58969, n58967, n58964, n58962, n58961,
         n58959, n58956, n58954, n58953, n58951, n58948, n58946, n58945,
         n58943, n58940, n58938, n58937, n58935, n58932, n58930, n58929,
         n58927, n58924, n58922, n58921, n58919, n58916, n58914, n58913,
         n58912, n58911, n58910, n58909, n58908, n58907, n58906, n58905,
         n58903, n58900, n58898, n58897, n58895, n58892, n58890, n58889,
         n58887, n58884, n58882, n58881, n58879, n58876, n58874, n58873,
         n58871, n58868, n58866, n58865, n58863, n58860, n58858, n58857,
         n58855, n58852, n58850, n58849, n58847, n58844, n58842, n58841,
         n58839, n58836, n58834, n58833, n58831, n58828, n58826, n58825,
         n58823, n58820, n58818, n58817, n58815, n58812, n58810, n58809,
         n58808, n58807, n58806, n58805, n58803, n58800, n58798, n58797,
         n58796, n58795, n58794, n58793, n58791, n58788, n58786, n58785,
         n58783, n58780, n58778, n58777, n58775, n58772, n58770, n58769,
         n58767, n58764, n58762, n58761, n58759, n58756, n58754, n58753,
         n58752, n58751, n58750, n58749, n58747, n58744, n58742, n58741,
         n58739, n58736, n58734, n58733, n58731, n58728, n58726, n58725,
         n58724, n58723, n58722, n58721, n58719, n58716, n58714, n58713,
         n58711, n58708, n58706, n58705, n58704, n58703, n58702, n58701,
         n58699, n58696, n58694, n58693, n58691, n58688, n58686, n58685,
         n58683, n58680, n58678, n58677, n58675, n58672, n58670, n58669,
         n58668, n58667, n58666, n58665, n58663, n58660, n58658, n58653,
         n58652, n58651, n58650, n58649, n58648, n58647, n58646, n58645,
         n58643, n58640, n58638, n58637, n58635, n58632, n58630, n58629,
         n58628, n58627, n58626, n58625, n58624, n58623, n58622, n58621,
         n58620, n58619, n58618, n58617, n58615, n58612, n58610, n58609,
         n58608, n58607, n58606, n58605, n58603, n58600, n58598, n58597,
         n58596, n58595, n58594, n58593, n58591, n58588, n58586, n58585,
         n58584, n58583, n58582, n58581, n58580, n58579, n58578, n58577,
         n58575, n58572, n58570, n58561, n58559, n58556, n58554, n58553,
         n58551, n58548, n58546, n58545, n58543, n58540, n58538, n58537,
         n58536, n58535, n58534, n58533, n58531, n58528, n58526, n58525,
         n58523, n58520, n58518, n58517, n58515, n58512, n58510, n58509,
         n58507, n58504, n58502, n58501, n58499, n58496, n58494, n58493,
         n58491, n58488, n58486, n58485, n58483, n58480, n58478, n58477,
         n58475, n58472, n58470, n58469, n58467, n58464, n58462, n58461,
         n58459, n58456, n58454, n58453, n58451, n58448, n58446, n58445,
         n58443, n58440, n58438, n58437, n58435, n58432, n58430, n58429,
         n58427, n58424, n58422, n58421, n58419, n58416, n58414, n58413,
         n58411, n58408, n58406, n58405, n58403, n58400, n58398, n58397,
         n58395, n58392, n58390, n58389, n58387, n58384, n58382, n58381,
         n58379, n58376, n58374, n58373, n58371, n58368, n58366, n58365,
         n58363, n58360, n58358, n58357, n58355, n58352, n58350, n58349,
         n58347, n58344, n58342, n58341, n58339, n58336, n58334, n58333,
         n58331, n58328, n58326, n58325, n58323, n58320, n58318, n58317,
         n58315, n58312, n58310, n58309, n58307, n58304, n58302, n58301,
         n58299, n58296, n58294, n58293, n58291, n58288, n58286, n58285,
         n58283, n58280, n58278, n58277, n58275, n58272, n58270, n58269,
         n58267, n58264, n58262, n58261, n58259, n58256, n58254, n58253,
         n58251, n58248, n58246, n58245, n58243, n58240, n58238, n58237,
         n58235, n58232, n58230, n58229, n58227, n58224, n58222, n58221,
         n58219, n58216, n58214, n58213, n58211, n58208, n58206, n58205,
         n58203, n58200, n58198, n58197, n58195, n58192, n58190, n58189,
         n58187, n58184, n58182, n58181, n58179, n58176, n58174, n58173,
         n58171, n58168, n58166, n58165, n58163, n58160, n58158, n58157,
         n58155, n58152, n58150, n58149, n58147, n58144, n58142, n58141,
         n58139, n58136, n58134, n58133, n58131, n58128, n58126, n58125,
         n58123, n58120, n58118, n58117, n58115, n58112, n58110, n58109,
         n58107, n58104, n58102, n58101, n58099, n58096, n58094, n58093,
         n58091, n58088, n58086, n58085, n58083, n58080, n58078, n58077,
         n58075, n58072, n58070, n58069, n58067, n58064, n58062, n58061,
         n58059, n58056, n58054, n58053, n58051, n58048, n58046, n58045,
         n58043, n58040, n58038, n58037, n58035, n58032, n58030, n58029,
         n58027, n58024, n58022, n58021, n58019, n58016, n58014, n58013,
         n58011, n58008, n58006, n58005, n58003, n58000, n57998, n57997,
         n57995, n57992, n57990, n57989, n57987, n57984, n57982, n57981,
         n57979, n57976, n57974, n57973, n57971, n57968, n57966, n57965,
         n57963, n57960, n57958, n57957, n57955, n57952, n57950, n57949,
         n57947, n57944, n57942, n57941, n57939, n57936, n57934, n57933,
         n57931, n57928, n57926, n57925, n57923, n57920, n57918, n57917,
         n57915, n57912, n57910, n57909, n57907, n57904, n57902, n57901,
         n57899, n57896, n57894, n57893, n57891, n57888, n57886, n57885,
         n57883, n57880, n57878, n57877, n57875, n57872, n57870, n57869,
         n57867, n57864, n57862, n57861, n57859, n57856, n57854, n57853,
         n57851, n57848, n57846, n57845, n57843, n57840, n57838, n57837,
         n57835, n57832, n57830, n57829, n57827, n57824, n57822, n57821,
         n57820, n57819, n57818, n57817, n57815, n57812, n57810, n57809,
         n57807, n57804, n57802, n57801, n57799, n57796, n57794, n57793,
         n57791, n57788, n57786, n57785, n57783, n57780, n57778, n57773,
         n57771, n57768, n57766, n57765, n57763, n57760, n57758, n57757,
         n57755, n57752, n57750, n57749, n57747, n57744, n57742, n57741,
         n57739, n57736, n57734, n57733, n57732, n57731, n57730, n57729,
         n57727, n57724, n57722, n57721, n57719, n57716, n57714, n57713,
         n57711, n57708, n57706, n57705, n57703, n57700, n57698, n57697,
         n57695, n57692, n57690, n57689, n57687, n57684, n57682, n57681,
         n57680, n57679, n57678, n57677, n57675, n57672, n57670, n57669,
         n57667, n57664, n57662, n57661, n57659, n57656, n57654, n57653,
         n57651, n57648, n57646, n57645, n57643, n57640, n57638, n57637,
         n57635, n57632, n57630, n57629, n57627, n57624, n57622, n57621,
         n57619, n57616, n57614, n57613, n57612, n57611, n57610, n57609,
         n57607, n57604, n57602, n57601, n57599, n57596, n57594, n57593,
         n57591, n57588, n57586, n57585, n57583, n57580, n57578, n57577,
         n57575, n57572, n57570, n57569, n57567, n57564, n57562, n57561,
         n57559, n57556, n57554, n57553, n57552, n57551, n57550, n57549,
         n57547, n57544, n57542, n57541, n57539, n57536, n57534, n57533,
         n57531, n57528, n57526, n57525, n57523, n57520, n57518, n57517,
         n57515, n57512, n57510, n57509, n57508, n57507, n57506, n57505,
         n57503, n57500, n57498, n57497, n57495, n57492, n57490, n57489,
         n57488, n57487, n57486, n57485, n57483, n57480, n57478, n57477,
         n57475, n57472, n57470, n57469, n57467, n57464, n57462, n57461,
         n57459, n57456, n57454, n57453, n57451, n57448, n57446, n57445,
         n57443, n57440, n57438, n57437, n57435, n57432, n57430, n57429,
         n57428, n57427, n57426, n57425, n57424, n57423, n57422, n57421,
         n57419, n57416, n57414, n57413, n57412, n57411, n57410, n57409,
         n57407, n57404, n57402, n57401, n57399, n57396, n57394, n57393,
         n57391, n57388, n57386, n57385, n57383, n57380, n57378, n57377,
         n57376, n57375, n57374, n57373, n57371, n57368, n57366, n57365,
         n57363, n57360, n57358, n57357, n57355, n57352, n57350, n57349,
         n57347, n57344, n57342, n57341, n57339, n57336, n57334, n57333,
         n57331, n57328, n57326, n57325, n57323, n57320, n57318, n57317,
         n57316, n57315, n57314, n57313, n57311, n57308, n57306, n57305,
         n57303, n57300, n57298, n57297, n57296, n57295, n57294, n57293,
         n57291, n57288, n57286, n57285, n57283, n57280, n57278, n57277,
         n57275, n57272, n57270, n57269, n57267, n57264, n57262, n57261,
         n57259, n57256, n57254, n57253, n57251, n57248, n57246, n57245,
         n57243, n57240, n57238, n57237, n57235, n57232, n57230, n57229,
         n57228, n57227, n57226, n57225, n57223, n57220, n57218, n57217,
         n57215, n57212, n57210, n57209, n57208, n57207, n57206, n57205,
         n57203, n57200, n57198, n57197, n57195, n57192, n57190, n57189,
         n57187, n57184, n57182, n57181, n57179, n57176, n57174, n57173,
         n57171, n57168, n57166, n57165, n57163, n57160, n57158, n57157,
         n57156, n57155, n57154, n57153, n57152, n57151, n57150, n57149,
         n57147, n57144, n57142, n57141, n57139, n57136, n57134, n57133,
         n57131, n57128, n57126, n57125, n57123, n57120, n57118, n57117,
         n57115, n57112, n57110, n57109, n57107, n57104, n57102, n57101,
         n57099, n57096, n57094, n57093, n57091, n57088, n57086, n57085,
         n57083, n57080, n57078, n57077, n57075, n57072, n57070, n57069,
         n57067, n57064, n57062, n57061, n57059, n57056, n57054, n57053,
         n57051, n57048, n57046, n57045, n57043, n57040, n57038, n57037,
         n57035, n57032, n57030, n57029, n57027, n57024, n57022, n57021,
         n57020, n57019, n57018, n57017, n57016, n57015, n57014, n57013,
         n57011, n57008, n57006, n57005, n57003, n57000, n56998, n56997,
         n56995, n56992, n56990, n56989, n56987, n56984, n56982, n56981,
         n56979, n56976, n56974, n56973, n56971, n56968, n56966, n56965,
         n56963, n56960, n56958, n56957, n56955, n56952, n56950, n56949,
         n56947, n56944, n56942, n56941, n56939, n56936, n56934, n56933,
         n56931, n56928, n56926, n56925, n56923, n56920, n56918, n56917,
         n56916, n56915, n56914, n56913, n56911, n56908, n56906, n56905,
         n56904, n56903, n56902, n56901, n56899, n56896, n56894, n56893,
         n56891, n56888, n56886, n56885, n56883, n56880, n56878, n56877,
         n56875, n56872, n56870, n56869, n56867, n56864, n56862, n56861,
         n56860, n56859, n56858, n56857, n56855, n56852, n56850, n56849,
         n56847, n56844, n56842, n56841, n56839, n56836, n56834, n56833,
         n56832, n56831, n56830, n56829, n56827, n56824, n56822, n56821,
         n56819, n56816, n56814, n56813, n56812, n56811, n56810, n56809,
         n56807, n56804, n56802, n56801, n56799, n56796, n56794, n56793,
         n56791, n56788, n56786, n56785, n56783, n56780, n56778, n56777,
         n56776, n56775, n56774, n56773, n56771, n56768, n56766, n56761,
         n56760, n56759, n56758, n56757, n56756, n56755, n56754, n56753,
         n56751, n56748, n56746, n56745, n56743, n56740, n56738, n56737,
         n56736, n56735, n56734, n56733, n56732, n56731, n56730, n56729,
         n56728, n56727, n56726, n56725, n56723, n56720, n56718, n56717,
         n56716, n56715, n56714, n56713, n56711, n56708, n56706, n56705,
         n56704, n56703, n56702, n56701, n56699, n56696, n56694, n56693,
         n56692, n56691, n56690, n56689, n56688, n56687, n56686, n56685,
         n56683, n56680, n56678, n56669, n56667, n56664, n56662, n56661,
         n56659, n56656, n56654, n56653, n56651, n56648, n56646, n56645,
         n56644, n56643, n56642, n56641, n56639, n56636, n56634, n56633,
         n56631, n56628, n56626, n56625, n56623, n56620, n56618, n56617,
         n56615, n56612, n56610, n56609, n56607, n56604, n56602, n56601,
         n56599, n56596, n56594, n56593, n56591, n56588, n56586, n56585,
         n56583, n56580, n56578, n56577, n56575, n56572, n56570, n56569,
         n56567, n56564, n56562, n56561, n56559, n56556, n56554, n56395,
         n56539, n56538, n56536, n56288, n56291, n56534, n56287, n56286,
         n56285, n56284, n56254, n56253, n56252, n56251, n56270, n56269,
         n56250, n56268, n56267, n56266, n56265, n56264, n56263, n56262,
         n56261, n56260, n56259, n56249, n56258, n56257, n56256, n56255,
         n56248, n64216, n64220, n64217, n64218, n64219, n56246, n56491,
         n56271, n56487, n56489, n56488, n56530, n56529, n56528, n56527,
         n56526, n56525, n56523, n56522, n56521, n56520, n56519, n56518,
         n56517, n56516, n56515, n56514, n56513, n56512, n56511, n56510,
         n56509, n56508, n56507, n56506, n56505, n56504, n56244, n56245,
         n56417, n56415, n56380, n56412, n56386, n56392, n56391, n56390,
         n56389, n64464, n56535, n56290, n64212, n64211, n56468, n56553,
         n56436, n60454, n60458, n60546, n61558, n64124, n56579, n56581,
         n56582, n56584, n58471, n58473, n58474, n58476, n60363, n60365,
         n60366, n60368, n62255, n62257, n62258, n62260, n62351, n62353,
         n62354, n62356, n56779, n56781, n56782, n56784, n58671, n58673,
         n58674, n58676, n60563, n60565, n60566, n60568, n62451, n62453,
         n62454, n62456, n56895, n56897, n56898, n56900, n58787, n58789,
         n58790, n58792, n60679, n60681, n60682, n60684, n62570, n62571,
         n62572, n62573, n62691, n62693, n62694, n62696, n57135, n57137,
         n57138, n57140, n59027, n59029, n59030, n59032, n60919, n60921,
         n60922, n60924, n57247, n57249, n57250, n57252, n59139, n59141,
         n59142, n59144, n61031, n61033, n61034, n61036, n62923, n62925,
         n62926, n62928, n57367, n57369, n57370, n57372, n59259, n59261,
         n59262, n59264, n61151, n61153, n61154, n61156, n63035, n63037,
         n63038, n63040, n57479, n57481, n57482, n57484, n59371, n59373,
         n59374, n59376, n61263, n61265, n61266, n61268, n57595, n57597,
         n57598, n57600, n59487, n59489, n59490, n59492, n61379, n61381,
         n61382, n61384, n63271, n63273, n63274, n63276, n57715, n57717,
         n57718, n57720, n59607, n59609, n59610, n59612, n61499, n61501,
         n61502, n61504, n63391, n63393, n63394, n63396, n57831, n57833,
         n57834, n57836, n59723, n59725, n59726, n59728, n61615, n61617,
         n61618, n61620, n63507, n63509, n63510, n63512, n57959, n57961,
         n57962, n57964, n59851, n59853, n59854, n59856, n61743, n61745,
         n61746, n61748, n63635, n63637, n63638, n63640, n58087, n58089,
         n58090, n58092, n59979, n59981, n59982, n59984, n61871, n61873,
         n61874, n61876, n63763, n63765, n63766, n63768, n58215, n58217,
         n58218, n58220, n60107, n60109, n60110, n60112, n61999, n62001,
         n62002, n62004, n63891, n63893, n63894, n63896, n58343, n58345,
         n58346, n58348, n60235, n60237, n60238, n60240, n62127, n62129,
         n62130, n62132, n64019, n64021, n64022, n64024, n56611, n56613,
         n56614, n56616, n58503, n58505, n58506, n58508, n60395, n60397,
         n60398, n60400, n62375, n62377, n62378, n62380, n62483, n62485,
         n62486, n62488, n56919, n56921, n56922, n56924, n58811, n58813,
         n58814, n58816, n60703, n60705, n60706, n60708, n62595, n62597,
         n62598, n62600, n57039, n57041, n57042, n57044, n58931, n58933,
         n58934, n58936, n60823, n60825, n60826, n60828, n62723, n62725,
         n62726, n62728, n57159, n57161, n57162, n57164, n59051, n59053,
         n59054, n59056, n60943, n60945, n60946, n60948, n62835, n62837,
         n62838, n62840, n57279, n57281, n57282, n57284, n59171, n59173,
         n59174, n59176, n61063, n61065, n61066, n61068, n57395, n57397,
         n57398, n57400, n59287, n59289, n59290, n59292, n61179, n61181,
         n61182, n61184, n63175, n63177, n63178, n63180, n57623, n57625,
         n57626, n57628, n59515, n59517, n59518, n59520, n61407, n61409,
         n61410, n61412, n63299, n63301, n63302, n63304, n57743, n57745,
         n57746, n57748, n59635, n59637, n59638, n59640, n61527, n61529,
         n61530, n61532, n63419, n63421, n63422, n63424, n57863, n57865,
         n57866, n57868, n59755, n59757, n59758, n59760, n61647, n61649,
         n61650, n61652, n63539, n63541, n63542, n63544, n57991, n57993,
         n57994, n57996, n59883, n59885, n59886, n59888, n61775, n61777,
         n61778, n61780, n63667, n63669, n63670, n63672, n58119, n58121,
         n58122, n58124, n60011, n60013, n60014, n60016, n61903, n61905,
         n61906, n61908, n63795, n63797, n63798, n63800, n58247, n58249,
         n58250, n58252, n60139, n60141, n60142, n60144, n62031, n62033,
         n62034, n62036, n63923, n63925, n63926, n63928, n58375, n58377,
         n58378, n58380, n60267, n60269, n60270, n60272, n62159, n62161,
         n62162, n62164, n64051, n64053, n64054, n64056, n62307, n62309,
         n62310, n62312, n62403, n62405, n62406, n62408, n56835, n56837,
         n56838, n56840, n58727, n58729, n58730, n58732, n60619, n60621,
         n60622, n60624, n62511, n62513, n62514, n62516, n56951, n56953,
         n56954, n56956, n58843, n58845, n58846, n58848, n60735, n60737,
         n60738, n60740, n62627, n62629, n62630, n62632, n57071, n57073,
         n57074, n57076, n58963, n58965, n58966, n58968, n60855, n60857,
         n60858, n60860, n62747, n62749, n62750, n62752, n57191, n57193,
         n57194, n57196, n59083, n59085, n59086, n59088, n60975, n60977,
         n60978, n60980, n62867, n62869, n62870, n62872, n57307, n57309,
         n57310, n57312, n59199, n59201, n59202, n59204, n61091, n61093,
         n61094, n61096, n62983, n62985, n62986, n62988, n63091, n63093,
         n63094, n63096, n57535, n57537, n57538, n57540, n59427, n59429,
         n59430, n59432, n61319, n61321, n61322, n61324, n63207, n63209,
         n63210, n63212, n57655, n57657, n57658, n57660, n59547, n59549,
         n59550, n59552, n61439, n61441, n61442, n61444, n63331, n63333,
         n63334, n63336, n57774, n57775, n57776, n57777, n59666, n59667,
         n59668, n59669, n61559, n61560, n61561, n63450, n63451, n63452,
         n63453, n57895, n57897, n57898, n57900, n59787, n59789, n59790,
         n59792, n61679, n61681, n61682, n61684, n63571, n63573, n63574,
         n63576, n58023, n58025, n58026, n58028, n59915, n59917, n59918,
         n59920, n61807, n61809, n61810, n61812, n63699, n63701, n63702,
         n63704, n58151, n58153, n58154, n58156, n60043, n60045, n60046,
         n60048, n61935, n61937, n61938, n61940, n63827, n63829, n63830,
         n63832, n58279, n58281, n58282, n58284, n60171, n60173, n60174,
         n60176, n62063, n62065, n62066, n62068, n63955, n63957, n63958,
         n63960, n58407, n58409, n58410, n58412, n60299, n60301, n60302,
         n60304, n62191, n62193, n62194, n62196, n64083, n64085, n64086,
         n64088, n56670, n56671, n56672, n56673, n58562, n58563, n58564,
         n58565, n60455, n60456, n60457, n62334, n62335, n62336, n62337,
         n62423, n62425, n62426, n62428, n56863, n56865, n56866, n56868,
         n58755, n58757, n58758, n58760, n60647, n60649, n60650, n60652,
         n62539, n62541, n62542, n62544, n56983, n56985, n56986, n56988,
         n58875, n58877, n58878, n58880, n60767, n60769, n60770, n60772,
         n62659, n62661, n62662, n62664, n57103, n57105, n57106, n57108,
         n58995, n58997, n58998, n59000, n60887, n60889, n60890, n60892,
         n62779, n62781, n62782, n62784, n57219, n57221, n57222, n57224,
         n59111, n59113, n59114, n59116, n61003, n61005, n61006, n61008,
         n57335, n57337, n57338, n57340, n59227, n59229, n59230, n59232,
         n61119, n61121, n61122, n61124, n57447, n57449, n57450, n57452,
         n59339, n59341, n59342, n59344, n61231, n61233, n61234, n61236,
         n63123, n63125, n63126, n63128, n57563, n57565, n57566, n57568,
         n59455, n59457, n59458, n59460, n61347, n61349, n61350, n61352,
         n63239, n63241, n63242, n63244, n57683, n57685, n57686, n57688,
         n59575, n59577, n59578, n59580, n61467, n61469, n61470, n61472,
         n63359, n63361, n63362, n63364, n57803, n57805, n57806, n57808,
         n59695, n59697, n59698, n59700, n61587, n61589, n61590, n61592,
         n63479, n63481, n63482, n63484, n57927, n57929, n57930, n57932,
         n59819, n59821, n59822, n59824, n61711, n61713, n61714, n61716,
         n63603, n63605, n63606, n63608, n58055, n58057, n58058, n58060,
         n59947, n59949, n59950, n59952, n61839, n61841, n61842, n61844,
         n63731, n63733, n63734, n63736, n58183, n58185, n58186, n58188,
         n60075, n60077, n60078, n60080, n61967, n61969, n61970, n61972,
         n63859, n63861, n63862, n63864, n58311, n58313, n58314, n58316,
         n60203, n60205, n60206, n60208, n62095, n62097, n62098, n62100,
         n63987, n63989, n63990, n63992, n58439, n58441, n58442, n58444,
         n60331, n60333, n60334, n60336, n62223, n62225, n62226, n62228,
         n64115, n64117, n64118, n64120, n56571, n56573, n56574, n56576,
         n58463, n58465, n58466, n58468, n60355, n60357, n60358, n60360,
         n62247, n62249, n62250, n62252, n62443, n62445, n62446, n62448,
         n56887, n56889, n56890, n56892, n58779, n58781, n58782, n58784,
         n60671, n60673, n60674, n60676, n62563, n62565, n62566, n62568,
         n57007, n57009, n57010, n57012, n58899, n58901, n58902, n58904,
         n60791, n60793, n60794, n60796, n62683, n62685, n62686, n62688,
         n57127, n57129, n57130, n57132, n59019, n59021, n59022, n59024,
         n60911, n60913, n60914, n60916, n62799, n62801, n62802, n62804,
         n57239, n57241, n57242, n57244, n59131, n59133, n59134, n59136,
         n61023, n61025, n61026, n61028, n62915, n62917, n62918, n62920,
         n57359, n57361, n57362, n57364, n59251, n59253, n59254, n59256,
         n61143, n61145, n61146, n61148, n63027, n63029, n63030, n63032,
         n57471, n57473, n57474, n57476, n59363, n59365, n59366, n59368,
         n61255, n61257, n61258, n61260, n63143, n63145, n63146, n63148,
         n57587, n57589, n57590, n57592, n59479, n59481, n59482, n59484,
         n61371, n61373, n61374, n61376, n63263, n63265, n63266, n63268,
         n57707, n57709, n57710, n57712, n59599, n59601, n59602, n59604,
         n61491, n61493, n61494, n61496, n63383, n63385, n63386, n63388,
         n57823, n57825, n57826, n57828, n59715, n59717, n59718, n59720,
         n61607, n61609, n61610, n61612, n63499, n63501, n63502, n63504,
         n57951, n57953, n57954, n57956, n59843, n59845, n59846, n59848,
         n61735, n61737, n61738, n61740, n63627, n63629, n63630, n63632,
         n58079, n58081, n58082, n58084, n59971, n59973, n59974, n59976,
         n61863, n61865, n61866, n61868, n63755, n63757, n63758, n63760,
         n58207, n58209, n58210, n58212, n60099, n60101, n60102, n60104,
         n61991, n61993, n61994, n61996, n63883, n63885, n63886, n63888,
         n58335, n58337, n58338, n58340, n60227, n60229, n60230, n60232,
         n62119, n62121, n62122, n62124, n64011, n64013, n64014, n64016,
         n56603, n56605, n56606, n56608, n58495, n58497, n58498, n58500,
         n60387, n60389, n60390, n60392, n56707, n56709, n56710, n56712,
         n58599, n58601, n58602, n58604, n60491, n60493, n60494, n60496,
         n62370, n62371, n62372, n62373, n56803, n56805, n56806, n56808,
         n58695, n58697, n58698, n58700, n60587, n60589, n60590, n60592,
         n62475, n62477, n62478, n62480, n62587, n62589, n62590, n62592,
         n57031, n57033, n57034, n57036, n58923, n58925, n58926, n58928,
         n60815, n60817, n60818, n60820, n62715, n62717, n62718, n62720,
         n62827, n62829, n62830, n62832, n57271, n57273, n57274, n57276,
         n59163, n59165, n59166, n59168, n61055, n61057, n61058, n61060,
         n62947, n62949, n62950, n62952, n57387, n57389, n57390, n57392,
         n59279, n59281, n59282, n59284, n61171, n61173, n61174, n61176,
         n63059, n63061, n63062, n63064, n57499, n57501, n57502, n57504,
         n59391, n59393, n59394, n59396, n61283, n61285, n61286, n61288,
         n63167, n63169, n63170, n63172, n57615, n57617, n57618, n57620,
         n59507, n59509, n59510, n59512, n61399, n61401, n61402, n61404,
         n63291, n63293, n63294, n63296, n57735, n57737, n57738, n57740,
         n59627, n59629, n59630, n59632, n61519, n61521, n61522, n61524,
         n63411, n63413, n63414, n63416, n57855, n57857, n57858, n57860,
         n59747, n59749, n59750, n59752, n61639, n61641, n61642, n61644,
         n63531, n63533, n63534, n63536, n57983, n57985, n57986, n57988,
         n59875, n59877, n59878, n59880, n61767, n61769, n61770, n61772,
         n63659, n63661, n63662, n63664, n58111, n58113, n58114, n58116,
         n60003, n60005, n60006, n60008, n61895, n61897, n61898, n61900,
         n63787, n63789, n63790, n63792, n58239, n58241, n58242, n58244,
         n60131, n60133, n60134, n60136, n62023, n62025, n62026, n62028,
         n63915, n63917, n63918, n63920, n58367, n58369, n58370, n58372,
         n60259, n60261, n60262, n60264, n62151, n62153, n62154, n62156,
         n64043, n64045, n64046, n64048, n56635, n56637, n56638, n56640,
         n58527, n58529, n58530, n58532, n60419, n60421, n60422, n60424,
         n62395, n62397, n62398, n62400, n62503, n62505, n62506, n62508,
         n56943, n56945, n56946, n56948, n58835, n58837, n58838, n58840,
         n60727, n60729, n60730, n60732, n62619, n62621, n62622, n62624,
         n57063, n57065, n57066, n57068, n58955, n58957, n58958, n58960,
         n60847, n60849, n60850, n60852, n62739, n62741, n62742, n62744,
         n57183, n57185, n57186, n57188, n59075, n59077, n59078, n59080,
         n60967, n60969, n60970, n60972, n62859, n62861, n62862, n62864,
         n57299, n57301, n57302, n57304, n59191, n59193, n59194, n59196,
         n61083, n61085, n61086, n61088, n62975, n62977, n62978, n62980,
         n57415, n57417, n57418, n57420, n59307, n59309, n59310, n59312,
         n61199, n61201, n61202, n61204, n57527, n57529, n57530, n57532,
         n59419, n59421, n59422, n59424, n61311, n61313, n61314, n61316,
         n63199, n63201, n63202, n63204, n57647, n57649, n57650, n57652,
         n59539, n59541, n59542, n59544, n61431, n61433, n61434, n61436,
         n63323, n63325, n63326, n63328, n57767, n57769, n57770, n57772,
         n59659, n59661, n59662, n59664, n61551, n61553, n61554, n61556,
         n63443, n63445, n63446, n63448, n57887, n57889, n57890, n57892,
         n59779, n59781, n59782, n59784, n61671, n61673, n61674, n61676,
         n63563, n63565, n63566, n63568, n58015, n58017, n58018, n58020,
         n59907, n59909, n59910, n59912, n61799, n61801, n61802, n61804,
         n63691, n63693, n63694, n63696, n58143, n58145, n58146, n58148,
         n60035, n60037, n60038, n60040, n61927, n61929, n61930, n61932,
         n63819, n63821, n63822, n63824, n58271, n58273, n58274, n58276,
         n60163, n60165, n60166, n60168, n62055, n62057, n62058, n62060,
         n63947, n63949, n63950, n63952, n58399, n58401, n58402, n58404,
         n60291, n60293, n60294, n60296, n62183, n62185, n62186, n62188,
         n64075, n64077, n64078, n64080, n56663, n56665, n56666, n56668,
         n58555, n58557, n58558, n58560, n60447, n60449, n60450, n60452,
         n62531, n62533, n62534, n62536, n56975, n56977, n56978, n56980,
         n58867, n58869, n58870, n58872, n60759, n60761, n60762, n60764,
         n62651, n62653, n62654, n62656, n57095, n57097, n57098, n57100,
         n58987, n58989, n58990, n58992, n60879, n60881, n60882, n60884,
         n62771, n62773, n62774, n62776, n57211, n57213, n57214, n57216,
         n59103, n59105, n59106, n59108, n60995, n60997, n60998, n61000,
         n62887, n62889, n62890, n62892, n57327, n57329, n57330, n57332,
         n59219, n59221, n59222, n59224, n61111, n61113, n61114, n61116,
         n57439, n57441, n57442, n57444, n59331, n59333, n59334, n59336,
         n61223, n61225, n61226, n61228, n63115, n63117, n63118, n63120,
         n57555, n57557, n57558, n57560, n59447, n59449, n59450, n59452,
         n61339, n61341, n61342, n61344, n63231, n63233, n63234, n63236,
         n57795, n57797, n57798, n57800, n59687, n59689, n59690, n59692,
         n61579, n61581, n61582, n61584, n63471, n63473, n63474, n63476,
         n57919, n57921, n57922, n57924, n59811, n59813, n59814, n59816,
         n61703, n61705, n61706, n61708, n63595, n63597, n63598, n63600,
         n58047, n58049, n58050, n58052, n59939, n59941, n59942, n59944,
         n61831, n61833, n61834, n61836, n63723, n63725, n63726, n63728,
         n58175, n58177, n58178, n58180, n60067, n60069, n60070, n60072,
         n61959, n61961, n61962, n61964, n63851, n63853, n63854, n63856,
         n58303, n58305, n58306, n58308, n60195, n60197, n60198, n60200,
         n62087, n62089, n62090, n62092, n63979, n63981, n63982, n63984,
         n58431, n58433, n58434, n58436, n60323, n60325, n60326, n60328,
         n62215, n62217, n62218, n62220, n64107, n64109, n64110, n64112,
         n56555, n56557, n56558, n56560, n58447, n58449, n58450, n58452,
         n60339, n60341, n60342, n60344, n62231, n62233, n62234, n62236,
         n56674, n56675, n56676, n56677, n58566, n58567, n58568, n58569,
         n60459, n60460, n60461, n62338, n62339, n62340, n62341, n56762,
         n56763, n56764, n56765, n58654, n58655, n58656, n58657, n60547,
         n60548, n60549, n62430, n62431, n62432, n62433, n56871, n56873,
         n56874, n56876, n58763, n58765, n58766, n58768, n60655, n60657,
         n60658, n60660, n62547, n62549, n62550, n62552, n56991, n56993,
         n56994, n56996, n58883, n58885, n58886, n58888, n60775, n60777,
         n60778, n60780, n62667, n62669, n62670, n62672, n57111, n57113,
         n57114, n57116, n59003, n59005, n59006, n59008, n60895, n60897,
         n60898, n60900, n62899, n62901, n62902, n62904, n57343, n57345,
         n57346, n57348, n59235, n59237, n59238, n59240, n61127, n61129,
         n61130, n61132, n63011, n63013, n63014, n63016, n57455, n57457,
         n57458, n57460, n59347, n59349, n59350, n59352, n61239, n61241,
         n61242, n61244, n57571, n57573, n57574, n57576, n59463, n59465,
         n59466, n59468, n61355, n61357, n61358, n61360, n63247, n63249,
         n63250, n63252, n57691, n57693, n57694, n57696, n59583, n59585,
         n59586, n59588, n61475, n61477, n61478, n61480, n63367, n63369,
         n63370, n63372, n57811, n57813, n57814, n57816, n59703, n59705,
         n59706, n59708, n61595, n61597, n61598, n61600, n63487, n63489,
         n63490, n63492, n57935, n57937, n57938, n57940, n59827, n59829,
         n59830, n59832, n61719, n61721, n61722, n61724, n63611, n63613,
         n63614, n63616, n58063, n58065, n58066, n58068, n59955, n59957,
         n59958, n59960, n61847, n61849, n61850, n61852, n63739, n63741,
         n63742, n63744, n58191, n58193, n58194, n58196, n60083, n60085,
         n60086, n60088, n61975, n61977, n61978, n61980, n63867, n63869,
         n63870, n63872, n58319, n58321, n58322, n58324, n60211, n60213,
         n60214, n60216, n62103, n62105, n62106, n62108, n63995, n63997,
         n63998, n64000, n56587, n56589, n56590, n56592, n58479, n58481,
         n58482, n58484, n60371, n60373, n60374, n60376, n62263, n62265,
         n62266, n62268, n56695, n56697, n56698, n56700, n58587, n58589,
         n58590, n58592, n60479, n60481, n60482, n60484, n62358, n62359,
         n62360, n62361, n56787, n56789, n56790, n56792, n58679, n58681,
         n58682, n58684, n60571, n60573, n60574, n60576, n62459, n62461,
         n62462, n62464, n62575, n62577, n62578, n62580, n62699, n62701,
         n62702, n62704, n57143, n57145, n57146, n57148, n59035, n59037,
         n59038, n59040, n60927, n60929, n60930, n60932, n62811, n62813,
         n62814, n62816, n57255, n57257, n57258, n57260, n59147, n59149,
         n59150, n59152, n61039, n61041, n61042, n61044, n62931, n62933,
         n62934, n62936, n63043, n63045, n63046, n63048, n57603, n57605,
         n57606, n57608, n59495, n59497, n59498, n59500, n61387, n61389,
         n61390, n61392, n63279, n63281, n63282, n63284, n57723, n57725,
         n57726, n57728, n59615, n59617, n59618, n59620, n61507, n61509,
         n61510, n61512, n63399, n63401, n63402, n63404, n57839, n57841,
         n57842, n57844, n59731, n59733, n59734, n59736, n61623, n61625,
         n61626, n61628, n63515, n63517, n63518, n63520, n57967, n57969,
         n57970, n57972, n59859, n59861, n59862, n59864, n61751, n61753,
         n61754, n61756, n63643, n63645, n63646, n63648, n58095, n58097,
         n58098, n58100, n59987, n59989, n59990, n59992, n61879, n61881,
         n61882, n61884, n63771, n63773, n63774, n63776, n58223, n58225,
         n58226, n58228, n60115, n60117, n60118, n60120, n62007, n62009,
         n62010, n62012, n63899, n63901, n63902, n63904, n58351, n58353,
         n58354, n58356, n60243, n60245, n60246, n60248, n62135, n62137,
         n62138, n62140, n64027, n64029, n64030, n64032, n56619, n56621,
         n56622, n56624, n58511, n58513, n58514, n58516, n60403, n60405,
         n60406, n60408, n62287, n62289, n62290, n62292, n56719, n56721,
         n56722, n56724, n58611, n58613, n58614, n58616, n60503, n60505,
         n60506, n60508, n56815, n56817, n56818, n56820, n58707, n58709,
         n58710, n58712, n60599, n60601, n60602, n60604, n56927, n56929,
         n56930, n56932, n58819, n58821, n58822, n58824, n60711, n60713,
         n60714, n60716, n62603, n62605, n62606, n62608, n57047, n57049,
         n57050, n57052, n58939, n58941, n58942, n58944, n60831, n60833,
         n60834, n60836, n57167, n57169, n57170, n57172, n59059, n59061,
         n59062, n59064, n60951, n60953, n60954, n60956, n62843, n62845,
         n62846, n62848, n57287, n57289, n57290, n57292, n59179, n59181,
         n59182, n59184, n61071, n61073, n61074, n61076, n62959, n62961,
         n62962, n62964, n57403, n57405, n57406, n57408, n59295, n59297,
         n59298, n59300, n61187, n61189, n61190, n61192, n63071, n63073,
         n63074, n63076, n57511, n57513, n57514, n57516, n59403, n59405,
         n59406, n59408, n61295, n61297, n61298, n61300, n63183, n63185,
         n63186, n63188, n57631, n57633, n57634, n57636, n59523, n59525,
         n59526, n59528, n61415, n61417, n61418, n61420, n63307, n63309,
         n63310, n63312, n57751, n57753, n57754, n57756, n59643, n59645,
         n59646, n59648, n61535, n61537, n61538, n61540, n63427, n63429,
         n63430, n63432, n57871, n57873, n57874, n57876, n59763, n59765,
         n59766, n59768, n61655, n61657, n61658, n61660, n63547, n63549,
         n63550, n63552, n57999, n58001, n58002, n58004, n59891, n59893,
         n59894, n59896, n61783, n61785, n61786, n61788, n63675, n63677,
         n63678, n63680, n58127, n58129, n58130, n58132, n60019, n60021,
         n60022, n60024, n61911, n61913, n61914, n61916, n63803, n63805,
         n63806, n63808, n58255, n58257, n58258, n58260, n60147, n60149,
         n60150, n60152, n62039, n62041, n62042, n62044, n63931, n63933,
         n63934, n63936, n58383, n58385, n58386, n58388, n60275, n60277,
         n60278, n60280, n62167, n62169, n62170, n62172, n64059, n64061,
         n64062, n64064, n56647, n56649, n56650, n56652, n58539, n58541,
         n58542, n58544, n60431, n60433, n60434, n60436, n62315, n62317,
         n62318, n62320, n56739, n56741, n56742, n56744, n58631, n58633,
         n58634, n58636, n60523, n60525, n60526, n60528, n56843, n56845,
         n56846, n56848, n58735, n58737, n58738, n58740, n60627, n60629,
         n60630, n60632, n62518, n62519, n62520, n62521, n56959, n56961,
         n56962, n56964, n58851, n58853, n58854, n58856, n60743, n60745,
         n60746, n60748, n62635, n62637, n62638, n62640, n57079, n57081,
         n57082, n57084, n58971, n58973, n58974, n58976, n60863, n60865,
         n60866, n60868, n62755, n62757, n62758, n62760, n57199, n57201,
         n57202, n57204, n59091, n59093, n59094, n59096, n60983, n60985,
         n60986, n60988, n63099, n63101, n63102, n63104, n57543, n57545,
         n57546, n57548, n59435, n59437, n59438, n59440, n61327, n61329,
         n61330, n61332, n63215, n63217, n63218, n63220, n57663, n57665,
         n57666, n57668, n59555, n59557, n59558, n59560, n61447, n61449,
         n61450, n61452, n63339, n63341, n63342, n63344, n57779, n57781,
         n57782, n57784, n59671, n59673, n59674, n59676, n61563, n61565,
         n61566, n61568, n63455, n63457, n63458, n63460, n57903, n57905,
         n57906, n57908, n59795, n59797, n59798, n59800, n61687, n61689,
         n61690, n61692, n63579, n63581, n63582, n63584, n58031, n58033,
         n58034, n58036, n59923, n59925, n59926, n59928, n61815, n61817,
         n61818, n61820, n63707, n63709, n63710, n63712, n58159, n58161,
         n58162, n58164, n60051, n60053, n60054, n60056, n61943, n61945,
         n61946, n61948, n63835, n63837, n63838, n63840, n58287, n58289,
         n58290, n58292, n60179, n60181, n60182, n60184, n62071, n62073,
         n62074, n62076, n63963, n63965, n63966, n63968, n58415, n58417,
         n58418, n58420, n60307, n60309, n60310, n60312, n62199, n62201,
         n62202, n62204, n64091, n64093, n64094, n64096, n56563, n56565,
         n56566, n56568, n58455, n58457, n58458, n58460, n60347, n60349,
         n60350, n60352, n62239, n62241, n62242, n62244, n56679, n56681,
         n56682, n56684, n58571, n58573, n58574, n58576, n60463, n60465,
         n60466, n60468, n62342, n62343, n62344, n62345, n56767, n56769,
         n56770, n56772, n58659, n58661, n58662, n58664, n60551, n60553,
         n60554, n60556, n62435, n62437, n62438, n62440, n56879, n56881,
         n56882, n56884, n58771, n58773, n58774, n58776, n60663, n60665,
         n60666, n60668, n62555, n62557, n62558, n62560, n56999, n57001,
         n57002, n57004, n58891, n58893, n58894, n58896, n60783, n60785,
         n60786, n60788, n62675, n62677, n62678, n62680, n57119, n57121,
         n57122, n57124, n59011, n59013, n59014, n59016, n60903, n60905,
         n60906, n60908, n62791, n62793, n62794, n62796, n57231, n57233,
         n57234, n57236, n59123, n59125, n59126, n59128, n61015, n61017,
         n61018, n61020, n62907, n62909, n62910, n62912, n57351, n57353,
         n57354, n57356, n59243, n59245, n59246, n59248, n61135, n61137,
         n61138, n61140, n63019, n63021, n63022, n63024, n57463, n57465,
         n57466, n57468, n59355, n59357, n59358, n59360, n61247, n61249,
         n61250, n61252, n63135, n63137, n63138, n63140, n57579, n57581,
         n57582, n57584, n59471, n59473, n59474, n59476, n61363, n61365,
         n61366, n61368, n63255, n63257, n63258, n63260, n57699, n57701,
         n57702, n57704, n59591, n59593, n59594, n59596, n61483, n61485,
         n61486, n61488, n63375, n63377, n63378, n63380, n57943, n57945,
         n57946, n57948, n59835, n59837, n59838, n59840, n61727, n61729,
         n61730, n61732, n63619, n63621, n63622, n63624, n58071, n58073,
         n58074, n58076, n59963, n59965, n59966, n59968, n61855, n61857,
         n61858, n61860, n63747, n63749, n63750, n63752, n58199, n58201,
         n58202, n58204, n60091, n60093, n60094, n60096, n61983, n61985,
         n61986, n61988, n63875, n63877, n63878, n63880, n58327, n58329,
         n58330, n58332, n60219, n60221, n60222, n60224, n62111, n62113,
         n62114, n62116, n64003, n64005, n64006, n64008, n56595, n56597,
         n56598, n56600, n58487, n58489, n58490, n58492, n60379, n60381,
         n60382, n60384, n62271, n62273, n62274, n62276, n62363, n62365,
         n62366, n62368, n56795, n56797, n56798, n56800, n58687, n58689,
         n58690, n58692, n60579, n60581, n60582, n60584, n62467, n62469,
         n62470, n62472, n56907, n56909, n56910, n56912, n58799, n58801,
         n58802, n58804, n60691, n60693, n60694, n60696, n57023, n57025,
         n57026, n57028, n58915, n58917, n58918, n58920, n60807, n60809,
         n60810, n60812, n62707, n62709, n62710, n62712, n62819, n62821,
         n62822, n62824, n57263, n57265, n57266, n57268, n59155, n59157,
         n59158, n59160, n61047, n61049, n61050, n61052, n62939, n62941,
         n62942, n62944, n57379, n57381, n57382, n57384, n59271, n59273,
         n59274, n59276, n61163, n61165, n61166, n61168, n63051, n63053,
         n63054, n63056, n57491, n57493, n57494, n57496, n59383, n59385,
         n59386, n59388, n61275, n61277, n61278, n61280, n63159, n63161,
         n63162, n63164, n57847, n57849, n57850, n57852, n59739, n59741,
         n59742, n59744, n61631, n61633, n61634, n61636, n63523, n63525,
         n63526, n63528, n57975, n57977, n57978, n57980, n59867, n59869,
         n59870, n59872, n61759, n61761, n61762, n61764, n63651, n63653,
         n63654, n63656, n58103, n58105, n58106, n58108, n59995, n59997,
         n59998, n60000, n61887, n61889, n61890, n61892, n63779, n63781,
         n63782, n63784, n58231, n58233, n58234, n58236, n60123, n60125,
         n60126, n60128, n62015, n62017, n62018, n62020, n63907, n63909,
         n63910, n63912, n58359, n58361, n58362, n58364, n60251, n60253,
         n60254, n60256, n62143, n62145, n62146, n62148, n64035, n64037,
         n64038, n64040, n56627, n56629, n56630, n56632, n58519, n58521,
         n58522, n58524, n60411, n60413, n60414, n60416, n62295, n62297,
         n62298, n62300, n62387, n62389, n62390, n62392, n56823, n56825,
         n56826, n56828, n58715, n58717, n58718, n58720, n60607, n60609,
         n60610, n60612, n62495, n62497, n62498, n62500, n56935, n56937,
         n56938, n56940, n58827, n58829, n58830, n58832, n60719, n60721,
         n60722, n60724, n62611, n62613, n62614, n62616, n57055, n57057,
         n57058, n57060, n58947, n58949, n58950, n58952, n60839, n60841,
         n60842, n60844, n57175, n57177, n57178, n57180, n59067, n59069,
         n59070, n59072, n60959, n60961, n60962, n60964, n62851, n62853,
         n62854, n62856, n62967, n62969, n62970, n62972, n63079, n63081,
         n63082, n63084, n57519, n57521, n57522, n57524, n59411, n59413,
         n59414, n59416, n61303, n61305, n61306, n61308, n63191, n63193,
         n63194, n63196, n57639, n57641, n57642, n57644, n59531, n59533,
         n59534, n59536, n61423, n61425, n61426, n61428, n63315, n63317,
         n63318, n63320, n57759, n57761, n57762, n57764, n59651, n59653,
         n59654, n59656, n61543, n61545, n61546, n61548, n63435, n63437,
         n63438, n63440, n57879, n57881, n57882, n57884, n59771, n59773,
         n59774, n59776, n61663, n61665, n61666, n61668, n63555, n63557,
         n63558, n63560, n58007, n58009, n58010, n58012, n59899, n59901,
         n59902, n59904, n61791, n61793, n61794, n61796, n63683, n63685,
         n63686, n63688, n58135, n58137, n58138, n58140, n60027, n60029,
         n60030, n60032, n61919, n61921, n61922, n61924, n63811, n63813,
         n63814, n63816, n58263, n58265, n58266, n58268, n60155, n60157,
         n60158, n60160, n62047, n62049, n62050, n62052, n63939, n63941,
         n63942, n63944, n58391, n58393, n58394, n58396, n60283, n60285,
         n60286, n60288, n62175, n62177, n62178, n62180, n64067, n64069,
         n64070, n64072, n56655, n56657, n56658, n56660, n58547, n58549,
         n58550, n58552, n60439, n60441, n60442, n60444, n62323, n62325,
         n62326, n62328, n56747, n56749, n56750, n56752, n58639, n58641,
         n58642, n58644, n60531, n60533, n60534, n60536, n56851, n56853,
         n56854, n56856, n58743, n58745, n58746, n58748, n60635, n60637,
         n60638, n60640, n62523, n62525, n62526, n62528, n56967, n56969,
         n56970, n56972, n58859, n58861, n58862, n58864, n60751, n60753,
         n60754, n60756, n62643, n62645, n62646, n62648, n57087, n57089,
         n57090, n57092, n58979, n58981, n58982, n58984, n60871, n60873,
         n60874, n60876, n62763, n62765, n62766, n62768, n62879, n62881,
         n62882, n62884, n57319, n57321, n57322, n57324, n59211, n59213,
         n59214, n59216, n61103, n61105, n61106, n61108, n62995, n62997,
         n62998, n63000, n57431, n57433, n57434, n57436, n59323, n59325,
         n59326, n59328, n61215, n61217, n61218, n61220, n63107, n63109,
         n63110, n63112, n63223, n63225, n63226, n63228, n57671, n57673,
         n57674, n57676, n59563, n59565, n59566, n59568, n61455, n61457,
         n61458, n61460, n63347, n63349, n63350, n63352, n57787, n57789,
         n57790, n57792, n59679, n59681, n59682, n59684, n61571, n61573,
         n61574, n61576, n63463, n63465, n63466, n63468, n57911, n57913,
         n57914, n57916, n59803, n59805, n59806, n59808, n61695, n61697,
         n61698, n61700, n63587, n63589, n63590, n63592, n58039, n58041,
         n58042, n58044, n59931, n59933, n59934, n59936, n61823, n61825,
         n61826, n61828, n63715, n63717, n63718, n63720, n58167, n58169,
         n58170, n58172, n60059, n60061, n60062, n60064, n61951, n61953,
         n61954, n61956, n63843, n63845, n63846, n63848, n58295, n58297,
         n58298, n58300, n60187, n60189, n60190, n60192, n62079, n62081,
         n62082, n62084, n63971, n63973, n63974, n63976, n58423, n58425,
         n58426, n58428, n60315, n60317, n60318, n60320, n62207, n62209,
         n62210, n62212, n64099, n64101, n64102, n64104, n56425, n56471,
         n56472, n56473, n56474, n56503, n56524, n56537, n56540, n56289,
         n56552, n56551, n56463, n56283, n56533, n56385, n64215, n23872,
         n23874, n23876, n23878, n23880, n23882, n23884, n23886, n23888,
         n23890, n23892, n23894, n23896, n23898, n23900, n23902, n23904,
         n23906, n23908, n23910, n23912, n23914, n23916, n23918, n23920,
         n23922, n23924, n23926, n23928, n23930, n23932, n23934, n23936,
         n23938, n23940, n23942, n23944, n23946, n23948, n23950, n23952,
         n23954, n23956, n23958, n23960, n23962, n23964, n23966, n23968,
         n23970, n23972, n23974, n23976, n23978, n23980, n23982, n23984,
         n23986, n23988, n23990, n23992, n23994, n23996, n23998, n24000,
         n24002, n24004, n24006, n24008, n24010, n24012, n24014, n24016,
         n24018, n24020, n24022, n24024, n24026, n24028, n24030, n24032,
         n24034, n24036, n24038, n24040, n24042, n24044, n24046, n24048,
         n24050, n24052, n24054, n24056, n24058, n24060, n24062, n24064,
         n24066, n24068, n24070, n24072, n24074, n24076, n24078, n24080,
         n24082, n24084, n24086, n24088, n24090, n24092, n24094, n24096,
         n24098, n24100, n24102, n24104, n24106, n24108, n24110, n24112,
         n24114, n24116, n24118, n24120, n24122, n24124, n24126, n24128,
         n24130, n24132, n24134, n24136, n24138, n24140, n24142, n24144,
         n24146, n24148, n24150, n24152, n24154, n24156, n24158, n24160,
         n24162, n24164, n24166, n24168, n24170, n24172, n24174, n24176,
         n24178, n24180, n24182, n24184, n24186, n24188, n24190, n24192,
         n24194, n24196, n24198, n24200, n24202, n24204, n24206, n24208,
         n24210, n24212, n24214, n24216, n24218, n24220, n24222, n24224,
         n24226, n24228, n24230, n24232, n24234, n24236, n24238, n24240,
         n24242, n24244, n24246, n24248, n24250, n24252, n24254, n24256,
         n24258, n24260, n24262, n24264, n24266, n24268, n24270, n24272,
         n24274, n24276, n24278, n24280, n24282, n24284, n24286, n24288,
         n24290, n24292, n24294, n24296, n24298, n24300, n24302, n24304,
         n24306, n24308, n24310, n24312, n24314, n24316, n24318, n24320,
         n24322, n24324, n24326, n24328, n24330, n24332, n24334, n24336,
         n24338, n24340, n24342, n24344, n24346, n24348, n24350, n24352,
         n24354, n24356, n24358, n24360, n24362, n24364, n24366, n24368,
         n24370, n24372, n24374, n24376, n24378, n24380, n24382, n24384,
         n24386, n24388, n24390, n24392, n24394, n24396, n24398, n24400,
         n24402, n24404, n24406, n24408, n24410, n24412, n24414, n24416,
         n24418, n24420, n24422, n24424, n24426, n24428, n24430, n24432,
         n24434, n24436, n24438, n24440, n24442, n24444, n24446, n24448,
         n24450, n24452, n24454, n24456, n24458, n24460, n24462, n24464,
         n24466, n24468, n24470, n24472, n24474, n24476, n24478, n24480,
         n24482, n24484, n24486, n24488, n24490, n24492, n24494, n24496,
         n24498, n24500, n24502, n24504, n24506, n24508, n24510, n24512,
         n24514, n24516, n24518, n24520, n24522, n24524, n24526, n24528,
         n24530, n24532, n24534, n24536, n24538, n24540, n24542, n24544,
         n24546, n24548, n24550, n24552, n24554, n24556, n24558, n24560,
         n24562, n24564, n24566, n24568, n24570, n24572, n24574, n24576,
         n24578, n24580, n24582, n24584, n24586, n24588, n24590, n24592,
         n24594, n24596, n24598, n24600, n24602, n24604, n24606, n24608,
         n24610, n24612, n24614, n24616, n24618, n24620, n24622, n24624,
         n24626, n24628, n24630, n24632, n24634, n24636, n24638, n24640,
         n24642, n24644, n24646, n24648, n24650, n24652, n24654, n24656,
         n24658, n24660, n24662, n24664, n24666, n24668, n24670, n24672,
         n24674, n24676, n24678, n24680, n24682, n24684, n24686, n24688,
         n24690, n24692, n24694, n24696, n24698, n24700, n24702, n24704,
         n24706, n24708, n24710, n24712, n24714, n24716, n24718, n24720,
         n24722, n24724, n24726, n24728, n24730, n24732, n24734, n24736,
         n24738, n24740, n24742, n24744, n24746, n24748, n24750, n24752,
         n24754, n24756, n24758, n24760, n24762, n24764, n24766, n24768,
         n24770, n24772, n24774, n24776, n24778, n24780, n24782, n24784,
         n24786, n24788, n24790, n24792, n24794, n24796, n24798, n24800,
         n24802, n24804, n24806, n24808, n24810, n24812, n24814, n24816,
         n24818, n24820, n24822, n24824, n24826, n24828, n24830, n24832,
         n24834, n24836, n24838, n24840, n24842, n24844, n24846, n24848,
         n24850, n24852, n24854, n24856, n24858, n24860, n24862, n24864,
         n24866, n24868, n24870, n24872, n24874, n24876, n24878, n24880,
         n24882, n24884, n24886, n24888, n24890, n24892, n24894, n24896,
         n24898, n24900, n24902, n24904, n24906, n24908, n24910, n24912,
         n24914, n24916, n24918, n24920, n24922, n24924, n24926, n24928,
         n24930, n24932, n24934, n24936, n24938, n24940, n24942, n24944,
         n24946, n24948, n24950, n24952, n24954, n24956, n24958, n24960,
         n24962, n24964, n24966, n24968, n24970, n24972, n24974, n24976,
         n24978, n24980, n24982, n24984, n24986, n24988, n24990, n24992,
         n24994, n24996, n24998, n25000, n25002, n25004, n25006, n25008,
         n25010, n25012, n25014, n25016, n25018, n25020, n25022, n25024,
         n25026, n25028, n25030, n25032, n25034, n25036, n25038, n25040,
         n25042, n25044, n25046, n25048, n25050, n25052, n25054, n25056,
         n25058, n25060, n25062, n25064, n25066, n25068, n25070, n25072,
         n25074, n25076, n25078, n25080, n25082, n25084, n25086, n25088,
         n25090, n25092, n25094, n25096, n25098, n25100, n25102, n25104,
         n25106, n25108, n25110, n25112, n25114, n25116, n25118, n25120,
         n25122, n25124, n25126, n25128, n25130, n25132, n25134, n25136,
         n25138, n25140, n25142, n25144, n25146, n25148, n25150, n25152,
         n25154, n25156, n25158, n25160, n25162, n25164, n25166, n25168,
         n25170, n25172, n25174, n25176, n25178, n25180, n25182, n25184,
         n25186, n25188, n25190, n25192, n25194, n25196, n25198, n25200,
         n25202, n25204, n25206, n25208, n25210, n25212, n25214, n25216,
         n25218, n25220, n25222, n25224, n25226, n25228, n25230, n25232,
         n25234, n25236, n25238, n25240, n25242, n25244, n25246, n25248,
         n25250, n25252, n25254, n25256, n25258, n25260, n25262, n25264,
         n25266, n25268, n25270, n25272, n25274, n25276, n25278, n25280,
         n25282, n25284, n25286, n25288, n25290, n25292, n25294, n25296,
         n25298, n25300, n25302, n25304, n25306, n25308, n25310, n25312,
         n25314, n25316, n25318, n25320, n25322, n25324, n25326, n25328,
         n25330, n25332, n25334, n25336, n25338, n25340, n25342, n25344,
         n25346, n25348, n25350, n25352, n25354, n25356, n25358, n25360,
         n25362, n25364, n25366, n25368, n25370, n25372, n25374, n25376,
         n25378, n25380, n25382, n25384, n25386, n25388, n25390, n25392,
         n25394, n25396, n25398, n25400, n25402, n25404, n25406, n25408,
         n25410, n25412, n25414, n25416, n25418, n25420, n25422, n25424,
         n25426, n25428, n25430, n25432, n25434, n25436, n25438, n25440,
         n25442, n25444, n25446, n25448, n25450, n25452, n25454, n25456,
         n25458, n25460, n25462, n25464, n25466, n25468, n25470, n25472,
         n25474, n25476, n25478, n25480, n25482, n25484, n25486, n25488,
         n25490, n25492, n25494, n25496, n25498, n25500, n25502, n25504,
         n25506, n25508, n25510, n25512, n25514, n25516, n25518, n25520,
         n25522, n25524, n25526, n25528, n25530, n25532, n25534, n25536,
         n25538, n25540, n25542, n25544, n25546, n25548, n25550, n25552,
         n25554, n25556, n25558, n25560, n25562, n25564, n25566, n25568,
         n25570, n25572, n25574, n25576, n25578, n25580, n25582, n25584,
         n25586, n25588, n25590, n25592, n25594, n25596, n25598, n25600,
         n25602, n25604, n25606, n25608, n25610, n25612, n25614, n25616,
         n25618, n25620, n25622, n25624, n25626, n25628, n25630, n25632,
         n25634, n25636, n25638, n25640, n25642, n25644, n25646, n25648,
         n25650, n25652, n25654, n25656, n25658, n25660, n25662, n25664,
         n25666, n25668, n25670, n25672, n25674, n25676, n25678, n25680,
         n25682, n25684, n25686, n25688, n25690, n25692, n25694, n25696,
         n25698, n25700, n25702, n25704, n25706, n25708, n25710, n25712,
         n25714, n25716, n25718, n25720, n25722, n25724, n25726, n25728,
         n25730, n25732, n25734, n25736, n25738, n25740, n25742, n25744,
         n25746, n25748, n25750, n25752, n25754, n25756, n25758, n25760,
         n25762, n25764, n25766, n25768, n25770, n25772, n25774, n25776,
         n25778, n25780, n25782, n25784, n25786, n25788, n25790, n25792,
         n25794, n25796, n25798, n25800, n25802, n25804, n25806, n25808,
         n25810, n25812, n25814, n25816, n25818, n25820, n25822, n25824,
         n25826, n25828, n25830, n25832, n25834, n25836, n25838, n25840,
         n25842, n25844, n25846, n25848, n25850, n25852, n25854, n25856,
         n25858, n25860, n25862, n25864, n25866, n25868, n25870, n25872,
         n25874, n25876, n25878, n25880, n25882, n25884, n25886, n25888,
         n25890, n25892, n25894, n25896, n25898, n25900, n25902, n25904,
         n25906, n25908, n25910, n25912, n25914, n25916, n25918, n25920,
         n25922, n25924, n25926, n25928, n25930, n25932, n25934, n25936,
         n25938, n25940, n25942, n25944, n25946, n25948, n25950, n25952,
         n25954, n25956, n25958, n25960, n25962, n25964, n25966, n25968,
         n25970, n25972, n25974, n25976, n25978, n25980, n25982, n25984,
         n25986, n25988, n25990, n25992, n25994, n25996, n25998, n26000,
         n26002, n26004, n26006, n26008, n26010, n26012, n26014, n26016,
         n26018, n26020, n26022, n26024, n26026, n26028, n26030, n26032,
         n26034, n26036, n26038, n26040, n26042, n26044, n26046, n26048,
         n26050, n26052, n26054, n26056, n26058, n26060, n26062, n26064,
         n26066, n26068, n26070, n26072, n26074, n26076, n26078, n26080,
         n26082, n26084, n26086, n26088, n26090, n26092, n26094, n26096,
         n26098, n26100, n26102, n26104, n26106, n26108, n26110, n26112,
         n26114, n26116, n26118, n26120, n26122, n26124, n26126, n26128,
         n26130, n26132, n26134, n26136, n26138, n26140, n26142, n26144,
         n26146, n26148, n26150, n26152, n26154, n26156, n26158, n26160,
         n26162, n26164, n26166, n26168, n26170, n26172, n26174, n26176,
         n26178, n26180, n26182, n26184, n26186, n26188, n26190, n26192,
         n26194, n26196, n26198, n26200, n26202, n26204, n26206, n26208,
         n26210, n26212, n26214, n26216, n26218, n26220, n26222, n26224,
         n26226, n26228, n26230, n26232, n26234, n26236, n26238, n26240,
         n26242, n26244, n26246, n26248, n26250, n26252, n26254, n26256,
         n26258, n26260, n26262, n26264, n26266, n26268, n26270, n26272,
         n26274, n26276, n26278, n26280, n26282, n26284, n26286, n26288,
         n26290, n26292, n26294, n26296, n26298, n26300, n26302, n26304,
         n26306, n26308, n26310, n26312, n26314, n26316, n26318, n26320,
         n26322, n26324, n26326, n26328, n26330, n26332, n26334, n26336,
         n26338, n26340, n26342, n26344, n26346, n26348, n26350, n26352,
         n26354, n26356, n26358, n26360, n26362, n26364, n26366, n26368,
         n26370, n26372, n26374, n26376, n26378, n26380, n26382, n26384,
         n26386, n26388, n26390, n26392, n26394, n26396, n26398, n26400,
         n26402, n26404, n26406, n26408, n26410, n26412, n26414, n26416,
         n26418, n26420, n26422, n26424, n26426, n26428, n26430, n26432,
         n26434, n26436, n26438, n26440, n26442, n26444, n26446, n26448,
         n26450, n26452, n26454, n26456, n26458, n26460, n26462, n26464,
         n26466, n26468, n26470, n26472, n26474, n26476, n26478, n26480,
         n26482, n26484, n26486, n26488, n26490, n26492, n26494, n26496,
         n26498, n26500, n26502, n26504, n26506, n26508, n26510, n26512,
         n26514, n26516, n26518, n26520, n26522, n26524, n26526, n26528,
         n26530, n26532, n26534, n26536, n26538, n26540, n26542, n26544,
         n26546, n26548, n26550, n26552, n26554, n26556, n26558, n26560,
         n26562, n26564, n26566, n26568, n26570, n26572, n26574, n26576,
         n26578, n26580, n26582, n26584, n26586, n26588, n26590, n26592,
         n26594, n26596, n26598, n26600, n26602, n26604, n26606, n26608,
         n26610, n26612, n26614, n26616, n26618, n26620, n26622, n26624,
         n26626, n26628, n26630, n26632, n26634, n26636, n26638, n26640,
         n26642, n26644, n26646, n26648, n26650, n26652, n26654, n26656,
         n26658, n26660, n26662, n26664, n26666, n26668, n26670, n26672,
         n26674, n26676, n26678, n26680, n26682, n26684, n26686, n26688,
         n26690, n26692, n26694, n26696, n26698, n26700, n26702, n26704,
         n26706, n26708, n26710, n26712, n26714, n26716, n26718, n26720,
         n26722, n26724, n26726, n26728, n26730, n26732, n26734, n26736,
         n26738, n26740, n26742, n26744, n26746, n26748, n26750, n26752,
         n26754, n26756, n26758, n26760, n26762, n26764, n26766, n26768,
         n26770, n26772, n26774, n26776, n26778, n26780, n26782, n26784,
         n26786, n26788, n26790, n26792, n26794, n26796, n26798, n26800,
         n26802, n26804, n26806, n26808, n26810, n26812, n26814, n26816,
         n26818, n26820, n26822, n26824, n26826, n26828, n26830, n26832,
         n26834, n26836, n26838, n26840, n26842, n26844, n26846, n26848,
         n26850, n26852, n26854, n26856, n26858, n26860, n26862, n26864,
         n26866, n26868, n26870, n26872, n26874, n26876, n26878, n26880,
         n26882, n26884, n26886, n26888, n26890, n26892, n26894, n26896,
         n26898, n26900, n26902, n26904, n26906, n26908, n26910, n26912,
         n26914, n26916, n26918, n26920, n26922, n26924, n26926, n26928,
         n26930, n26932, n26934, n26936, n26938, n26940, n26942, n26944,
         n26946, n26948, n26950, n26952, n26954, n26956, n26958, n26960,
         n26962, n26964, n26966, n26968, n26970, n26972, n26974, n26976,
         n26978, n26980, n26982, n26984, n26986, n26988, n26990, n26992,
         n26994, n26996, n26998, n27000, n27002, n27004, n27006, n27008,
         n27010, n27012, n27014, n27016, n27018, n27020, n27022, n27024,
         n27026, n27028, n27030, n27032, n27034, n27036, n27038, n27040,
         n27042, n27044, n27046, n27048, n27050, n27052, n27054, n27056,
         n27058, n27060, n27062, n27064, n27066, n27068, n27070, n27072,
         n27074, n27076, n27078, n27080, n27082, n27084, n27086, n27088,
         n27090, n27092, n27094, n27096, n27098, n27100, n27102, n27104,
         n27106, n27108, n27110, n27112, n27114, n27116, n27118, n27120,
         n27122, n27124, n27126, n27128, n27130, n27132, n27134, n27136,
         n27138, n27140, n27142, n27144, n27146, n27148, n27150, n27152,
         n27154, n27156, n27158, n27160, n27162, n27164, n27166, n27168,
         n27170, n27172, n27174, n27176, n27178, n27180, n27182, n27184,
         n27186, n27188, n27190, n27192, n27194, n27196, n27198, n27200,
         n27202, n27204, n27206, n27208, n27210, n27212, n27214, n27216,
         n27218, n27220, n27222, n27224, n27226, n27228, n27230, n27232,
         n27234, n27236, n27238, n27240, n27242, n27244, n27246, n27248,
         n27250, n27252, n27254, n27256, n27258, n27260, n27262, n27264,
         n27266, n27268, n27270, n27272, n27274, n27276, n27278, n27280,
         n27282, n27284, n27286, n27288, n27290, n27292, n27294, n27296,
         n27298, n27300, n27302, n27304, n27306, n27308, n27310, n27312,
         n27314, n27316, n27318, n27320, n27322, n27324, n27326, n27328,
         n27330, n27332, n27334, n27336, n27338, n27340, n27342, n27344,
         n27346, n27348, n27350, n27352, n27354, n27356, n27358, n27360,
         n27362, n27364, n27366, n27368, n27370, n27372, n27374, n27376,
         n27378, n27380, n27382, n27384, n27386, n27388, n27390, n27392,
         n27394, n27396, n27398, n27400, n27402, n27404, n27406, n27408,
         n27410, n27412, n27414, n27416, n27418, n27420, n27422, n27424,
         n27426, n27428, n27430, n27432, n27434, n27436, n27438, n27440,
         n27442, n27444, n27446, n27448, n27450, n27452, n27454, n27456,
         n27458, n27460, n27462, n27464, n27466, n27468, n27470, n27472,
         n27474, n27476, n27478, n27480, n27482, n27484, n27486, n27488,
         n27490, n27492, n27494, n27496, n27498, n27500, n27502, n27504,
         n27506, n27508, n27510, n27512, n27514, n27516, n27518, n27520,
         n27522, n27524, n27526, n27528, n27530, n27532, n27534, n27536,
         n27538, n27540, n27542, n27544, n27546, n27548, n27550, n27552,
         n27554, n27556, n27558, n27560, n27562, n27564, n27566, n27568,
         n27570, n27572, n27574, n27576, n27578, n27580, n27582, n27584,
         n27586, n27588, n27590, n27592, n27594, n27596, n27598, n27600,
         n27602, n27604, n27606, n27608, n27610, n27612, n27614, n27616,
         n27618, n27620, n27622, n27624, n27626, n27628, n27630, n27632,
         n27634, n27636, n27638, n27640, n27642, n27644, n27646, n27648,
         n27650, n27652, n27654, n27656, n27658, n27660, n27662, n27664,
         n27666, n27668, n27670, n27672, n27674, n27676, n27678, n27680,
         n27682, n27684, n27686, n27688, n27690, n27692, n27694, n27696,
         n27698, n27700, n27702, n27704, n27706, n27708, n27710, n27712,
         n27714, n27716, n27718, n27720, n27722, n27724, n27726, n27728,
         n27730, n27732, n27734, n27736, n27738, n27740, n27742, n27744,
         n27746, n27748, n27750, n27752, n27754, n27756, n27758, n27760,
         n27762, n27764, n27766, n27768, n27770, n27772, n27774, n27776,
         n27778, n27780, n27782, n27784, n27786, n27788, n27790, n27792,
         n27794, n27796, n27798, n27800, n27802, n27804, n27806, n27808,
         n27810, n27812, n27814, n27816, n27818, n27820, n27822, n27824,
         n27826, n27828, n27830, n27832, n27834, n27836, n27838, n27840,
         n27842, n27844, n27846, n27848, n27850, n27852, n27854, n27856,
         n27858, n27860, n27862, n27864, n27866, n27868, n27870, n27872,
         n27874, n27876, n27878, n27880, n27882, n27884, n27886, n27888,
         n27890, n27892, n27894, n27896, n27898, n27900, n27902, n27904,
         n27906, n27908, n27910, n27912, n27914, n27916, n27918, n27920,
         n27922, n27924, n27926, n27928, n27930, n27932, n27934, n27936,
         n27938, n27940, n27942, n27944, n27946, n27948, n27950, n27952,
         n27954, n27956, n27958, n27960, n27962, n27964, n27966, n27968,
         n27970, n27972, n27974, n27976, n27978, n27980, n27982, n27984,
         n27986, n27988, n27990, n27992, n27994, n27996, n27998, n28000,
         n28002, n28004, n28006, n28008, n28010, n28012, n28014, n28016,
         n28018, n28020, n28022, n28024, n28026, n28028, n28030, n28032,
         n28034, n28036, n28038, n28040, n28042, n28044, n28046, n28048,
         n28050, n28052, n28054, n28056, n28058, n28060, n28062, n28064,
         n28066, n28068, n28070, n28072, n28074, n28076, n28078, n28080,
         n28082, n28084, n28086, n28088, n28090, n28092, n28094, n28096,
         n28098, n28100, n28102, n28104, n28106, n28108, n28110, n28112,
         n28114, n28116, n28118, n28120, n28122, n28124, n28126, n28128,
         n28130, n28132, n28134, n28136, n28138, n28140, n28142, n28144,
         n28146, n28148, n28150, n28152, n28154, n28156, n28158, n28160,
         n28162, n28164, n28166, n28168, n28170, n28172, n28174, n28176,
         n28178, n28180, n28182, n28184, n28186, n28188, n28190, n28192,
         n28194, n28196, n28198, n28200, n28202, n28204, n28206, n28208,
         n28210, n28212, n28214, n28216, n28218, n28220, n28222, n28224,
         n28226, n28228, n28230, n28232, n28234, n28236, n28238, n28240,
         n28242, n28244, n28246, n28248, n28250, n28252, n28254, n28256,
         n28258, n28260, n28262, n28264, n28266, n28268, n28270, n28272,
         n28274, n28276, n28278, n28280, n28282, n28284, n28286, n28288,
         n28290, n28292, n28294, n28296, n28298, n28300, n28302, n28304,
         n28306, n28308, n28310, n28312, n28314, n28316, n28318, n28320,
         n28322, n28324, n28326, n28328, n28330, n28332, n28334, n28336,
         n28338, n28340, n28342, n28344, n28346, n28348, n28350, n28352,
         n28354, n28356, n28358, n28360, n28362, n28364, n28366, n28368,
         n28370, n28372, n28374, n28376, n28378, n28380, n28382, n28384,
         n28386, n28388, n28390, n28392, n28394, n28396, n28398, n28400,
         n28402, n28404, n28406, n28408, n28410, n28412, n28414, n28416,
         n28418, n28420, n28422, n28424, n28426, n28428, n28430, n28432,
         n28434, n28436, n28438, n28440, n28442, n28444, n28446, n28448,
         n28450, n28452, n28454, n28456, n28458, n28460, n28462, n28464,
         n28466, n28468, n28470, n28472, n28474, n28476, n28478, n28480,
         n28482, n28484, n28486, n28488, n28490, n28492, n28494, n28496,
         n28498, n28500, n28502, n28504, n28506, n28508, n28510, n28512,
         n28514, n28516, n28518, n28520, n28522, n28524, n28526, n28528,
         n28530, n28532, n28534, n28536, n28538, n28540, n28542, n28544,
         n28546, n28548, n28550, n28552, n28554, n28556, n28558, n28560,
         n28562, n28564, n28566, n28568, n28570, n28572, n28574, n28576,
         n28578, n28580, n28582, n28584, n28586, n28588, n28590, n28592,
         n28594, n28596, n28598, n28600, n28602, n28604, n28606, n28608,
         n28610, n28612, n28614, n28616, n28618, n28620, n28622, n28624,
         n28626, n28628, n28630, n28632, n28634, n28636, n28638, n28640,
         n28642, n28644, n28646, n28648, n28650, n28652, n28654, n28656,
         n28658, n28660, n28662, n28664, n28666, n28668, n28670, n28672,
         n28674, n28676, n28678, n28680, n28682, n28684, n28686, n28688,
         n28690, n28692, n28694, n28696, n28698, n28700, n28702, n28704,
         n28706, n28708, n28710, n28712, n28714, n28716, n28718, n28720,
         n28722, n28724, n28726, n28728, n28730, n28732, n28734, n28736,
         n28738, n28740, n28742, n28744, n28746, n28748, n28750, n28752,
         n28754, n28756, n28758, n28760, n28762, n28764, n28766, n28768,
         n28770, n28772, n28774, n28776, n28778, n28780, n28782, n28784,
         n28786, n28788, n28790, n28792, n28794, n28796, n28798, n28800,
         n28802, n28804, n28806, n28808, n28810, n28812, n28814, n28816,
         n28818, n28820, n28822, n28824, n28826, n28828, n28830, n28832,
         n28834, n28836, n28838, n28840, n28842, n28844, n28846, n28848,
         n28850, n28852, n28854, n28856, n28858, n28860, n28862, n28864,
         n28866, n28868, n28870, n28872, n28874, n28876, n28878, n28880,
         n28882, n28884, n28886, n28888, n28890, n28892, n28894, n28896,
         n28898, n28900, n28902, n28904, n28906, n28908, n28910, n28912,
         n28914, n28916, n28918, n28920, n28922, n28924, n28926, n28928,
         n28930, n28932, n28934, n28936, n28938, n28940, n28942, n28944,
         n28946, n28948, n28950, n28952, n28954, n28956, n28958, n28960,
         n28962, n28964, n28966, n28968, n28970, n28972, n28974, n28976,
         n28978, n28980, n28982, n28984, n28986, n28988, n28990, n28992,
         n28994, n28996, n28998, n29000, n29002, n29004, n29006, n29008,
         n29010, n29012, n29014, n29016, n29018, n29020, n29022, n29024,
         n29026, n29028, n29030, n29032, n29034, n29036, n29038, n29040,
         n29042, n29044, n29046, n29048, n29050, n29052, n29054, n29056,
         n29058, n29060, n29062, n29064, n29066, n29068, n29070, n29072,
         n29074, n29076, n29078, n29080, n29082, n29084, n29086, n29088,
         n29090, n29092, n29094, n29096, n29098, n29100, n29102, n29104,
         n29106, n29108, n29110, n29112, n29114, n29116, n29118, n29120,
         n29122, n29124, n29126, n29128, n29130, n29132, n29134, n29136,
         n29138, n29140, n29142, n29144, n29146, n29148, n29150, n29152,
         n29154, n29156, n29158, n29160, n29162, n29164, n29166, n29168,
         n29170, n29172, n29174, n29176, n29178, n29180, n29182, n29184,
         n29186, n29188, n29190, n29192, n29194, n29196, n29198, n29200,
         n29202, n29204, n29206, n29208, n29210, n29212, n29214, n29216,
         n29218, n29220, n29222, n29224, n29226, n29228, n29230, n29232,
         n29234, n29236, n29238, n29240, n29242, n29244, n29246, n29248,
         n29250, n29252, n29254, n29256, n29258, n29260, n29262, n29264,
         n29266, n29268, n29270, n29272, n29274, n29276, n29278, n29280,
         n29282, n29284, n29286, n29288, n29290, n29292, n29294, n29296,
         n29298, n29300, n29302, n29304, n29306, n29308, n29310, n29312,
         n29314, n29316, n29318, n29320, n29322, n29324, n29326, n29328,
         n29330, n29332, n29334, n29336, n29338, n29340, n29342, n29344,
         n29346, n29348, n29350, n29352, n29354, n29356, n29358, n29360,
         n29362, n29364, n29366, n29368, n29370, n29372, n29374, n29376,
         n29378, n29380, n29382, n29384, n29386, n29388, n29390, n29392,
         n29394, n29396, n29398, n29400, n29402, n29404, n29406, n29408,
         n29410, n29412, n29414, n29416, n29418, n29420, n29422, n29424,
         n29426, n29428, n29430, n29432, n29434, n29436, n29438, n29440,
         n29442, n29444, n29446, n29448, n29450, n29452, n29454, n29456,
         n29458, n29460, n29462, n29464, n29466, n29468, n29470, n29472,
         n29474, n29476, n29478, n29480, n29482, n29484, n29486, n29488,
         n29490, n29492, n29494, n29496, n29498, n29500, n29502, n29504,
         n29506, n29508, n29510, n29512, n29514, n29516, n29518, n29520,
         n29522, n29524, n29526, n29528, n29530, n29532, n29534, n29536,
         n29538, n29540, n29542, n29544, n29546, n29548, n29550, n29552,
         n29554, n29556, n29558, n29560, n29562, n29564, n29566, n29568,
         n29570, n29572, n29574, n29576, n29578, n29580, n29582, n29584,
         n29586, n29588, n29590, n29592, n29594, n29596, n29598, n29600,
         n29602, n29604, n29606, n29608, n29610, n29612, n29614, n29616,
         n29618, n29620, n29622, n29624, n29626, n29628, n29630, n29632,
         n29634, n29636, n29638, n29640, n29642, n29644, n29646, n29648,
         n29650, n29652, n29654, n29656, n29658, n29660, n29662, n29664,
         n29666, n29668, n29670, n29672, n29674, n29676, n29678, n29680,
         n29682, n29684, n29686, n29688, n29690, n29692, n29694, n29696,
         n29698, n29700, n29702, n29704, n29706, n29708, n29710, n29712,
         n29714, n29716, n29718, n29720, n29722, n29724, n29726, n29728,
         n29730, n29732, n29734, n29736, n29738, n29740, n29742, n29744,
         n29746, n29748, n29750, n29752, n29754, n29756, n29758, n29760,
         n29762, n29764, n29766, n29768, n29770, n29772, n29774, n29776,
         n29778, n29780, n29782, n29784, n29786, n29788, n29790, n29792,
         n29794, n29796, n29798, n29800, n29802, n29804, n29806, n29808,
         n29810, n29812, n29814, n29816, n29818, n29820, n29822, n29824,
         n29826, n29828, n29830, n29832, n29834, n29836, n29838, n29840,
         n29842, n29844, n29846, n29848, n29850, n29852, n29854, n29856,
         n29858, n29860, n29862, n29864, n29866, n29868, n29870, n29872,
         n29874, n29876, n29878, n29880, n29882, n29884, n29886, n29888,
         n29890, n29892, n29894, n29896, n29898, n29900, n29902, n29904,
         n29906, n29908, n29910, n29912, n29914, n29916, n29918, n29920,
         n29922, n29924, n29926, n29928, n29930, n29932, n29934, n29936,
         n29938, n29940, n29942, n29944, n29946, n29948, n29950, n29952,
         n29954, n29956, n29958, n29960, n29962, n29964, n29966, n29968,
         n29970, n29972, n29974, n29976, n29978, n29980, n29982, n29984,
         n29986, n29988, n29990, n29992, n29994, n29996, n29998, n30000,
         n30002, n30004, n30006, n30008, n30010, n30012, n30014, n30016,
         n30018, n30020, n30022, n30024, n30026, n30028, n30030, n30032,
         n30034, n30036, n30038, n30040, n30042, n30044, n30046, n30048,
         n30050, n30052, n30054, n30056, n30058, n30060, n30062, n30064,
         n30066, n30068, n30070, n30072, n30074, n30076, n30078, n30080,
         n30082, n30084, n30086, n30088, n30090, n30092, n30094, n30096,
         n30098, n30100, n30102, n30104, n30106, n30108, n30110, n30112,
         n30114, n30116, n30118, n30120, n30122, n30124, n30126, n30128,
         n30130, n30132, n30134, n30136, n30138, n30140, n30142, n30144,
         n30146, n30148, n30150, n30152, n30154, n30156, n30158, n30160,
         n30162, n30164, n30166, n30168, n30170, n30172, n30174, n30176,
         n30178, n30180, n30182, n30184, n30186, n30188, n30190, n30192,
         n30194, n30196, n30198, n30200, n30202, n30204, n30206, n30208,
         n30210, n30212, n30214, n30216, n30218, n30220, n30222, n30224,
         n30226, n30228, n30230, n30232, n30234, n30236, n30238, n30240,
         n30242, n30244, n30246, n30248, n30250, n30252, n30254, n30256,
         n30258, n30260, n30262, n30264, n30266, n30268, n30270, n30272,
         n30274, n30276, n30278, n30280, n30282, n30284, n30286, n30288,
         n30290, n30292, n30294, n30296, n30298, n30300, n30302, n30304,
         n30306, n30308, n30310, n30312, n30314, n30316, n30318, n30320,
         n30322, n30324, n30326, n30328, n30330, n30332, n30334, n30336,
         n30338, n30340, n30342, n30344, n30346, n30348, n30350, n30352,
         n30354, n30356, n30358, n30360, n30362, n30364, n30366, n30368,
         n30370, n30372, n30374, n30376, n30378, n30380, n30382, n30384,
         n30386, n30388, n30390, n30392, n30394, n30396, n30398, n30400,
         n30402, n30404, n30406, n30408, n30410, n30412, n30414, n30416,
         n30418, n30420, n30422, n30424, n30426, n30428, n30430, n30432,
         n30434, n30436, n30438, n30440, n30442, n30444, n30446, n30448,
         n30450, n30452, n30454, n30456, n30458, n30460, n30462, n30464,
         n30466, n30468, n30470, n30472, n30474, n30476, n30478, n30480,
         n30482, n30484, n30486, n30488, n30490, n30492, n30494, n30496,
         n30498, n30500, n30502, n30504, n30506, n30508, n30510, n30512,
         n30514, n30516, n30518, n30520, n30522, n30524, n30526, n30528,
         n30530, n30532, n30534, n30536, n30538, n30540, n30542, n30544,
         n30546, n30548, n30550, n30552, n30554, n30556, n30558, n30560,
         n30562, n30564, n30566, n30568, n30570, n30572, n30574, n30576,
         n30578, n30580, n30582, n30584, n30586, n30588, n30590, n30592,
         n30594, n30596, n30598, n30600, n30602, n30604, n30606, n30608,
         n30610, n30612, n30614, n30616, n30618, n30620, n30622, n30624,
         n30626, n30628, n30630, n30632, n30634, n30636, n30638, n30640,
         n30642, n30644, n30646, n30648, n30650, n30652, n30654, n30656,
         n30658, n30660, n30662, n30664, n30666, n30668, n30670, n30672,
         n30674, n30676, n30678, n30680, n30682, n30684, n30686, n30688,
         n30690, n30692, n30694, n30696, n30698, n30700, n30702, n30704,
         n30706, n30708, n30710, n30712, n30714, n30716, n30718, n30720,
         n30722, n30724, n30726, n30728, n30730, n30732, n30734, n30736,
         n30738, n30740, n30742, n30744, n30746, n30748, n30750, n30752,
         n30754, n30756, n30758, n30760, n30762, n30764, n30766, n30768,
         n30770, n30772, n30774, n30776, n30778, n30780, n30782, n30784,
         n30786, n30788, n30790, n30792, n30794, n30796, n30798, n30800,
         n30802, n30804, n30806, n30808, n30810, n30812, n30814, n30816,
         n30818, n30820, n30822, n30824, n30826, n30828, n30830, n30832,
         n30834, n30836, n30838, n30840, n30842, n30844, n30846, n30848,
         n30850, n30852, n30854, n30856, n30858, n30860, n30862, n30864,
         n30866, n30868, n30870, n30872, n30874, n30876, n30878, n30880,
         n30882, n30884, n30886, n30888, n30890, n30892, n30894, n30896,
         n30898, n30900, n30902, n30904, n30906, n30908, n30910, n30912,
         n30914, n30916, n30918, n30920, n30922, n30924, n30926, n30928,
         n30930, n30932, n30934, n30936, n30938, n30940, n30942, n30944,
         n30946, n30948, n30950, n30952, n30954, n30956, n30958, n30960,
         n30962, n30964, n30966, n30968, n30970, n30972, n30974, n30976,
         n30978, n30980, n30982, n30984, n30986, n30988, n30990, n30992,
         n30994, n30996, n30998, n31000, n31002, n31004, n31006, n31008,
         n31010, n31012, n31014, n31016, n31018, n31020, n31022, n31024,
         n31026, n31028, n31030, n31032, n31034, n31036, n31038, n31040,
         n31042, n31044, n31046, n31048, n31050, n31052, n31054, n31056,
         n31058, n31060, n31062, n31064, n31066, n31068, n31070, n31072,
         n31074, n31076, n31078, n31080, n31082, n31084, n31086, n31088,
         n31090, n31092, n31094, n31096, n31098, n31100, n31102, n31104,
         n31106, n31108, n31110, n31112, n31114, n31116, n31118, n31120,
         n31122, n31124, n31126, n31128, n31130, n31132, n31134, n31136,
         n31138, n31140, n31142, n31144, n31146, n31148, n31150, n31152,
         n31154, n31156, n31158, n31160, n31162, n31164, n31166, n31168,
         n31170, n31172, n31174, n31176, n31178, n31180, n31182, n31184,
         n31186, n31188, n31190, n31192, n31194, n31196, n31198, n31200,
         n31202, n31204, n31206, n31208, n31210, n31212, n31214, n31216,
         n31218, n31220, n31222, n31224, n31226, n31228, n31230, n31232,
         n31234, n31236, n31238, n31240, n31242, n31244, n31246, n31248,
         n31250, n31252, n31254, n31256, n31258, n31260, n31262, n31264,
         n31266, n31268, n31270, n31272, n31274, n31276, n31278, n31280,
         n31282, n31284, n31286, n31288, n31290, n31292, n31294, n31296,
         n31298, n31300, n31302, n31304, n31306, n31308, n31310, n31312,
         n31314, n31316, n31318, n31320, n31322, n31324, n31326, n31328,
         n31330, n31332, n31334, n31336, n31338, n31341, n31343, n31345,
         n31347, n31349, n31351, n31353, n31356, n31358, n31360, n31362,
         n31364, n31367, n31369, n31371, n31373, n31375, n31378, n31380,
         n31382, n31384, n31386, n31389, n31391, n31393, n31395, n31397,
         n31399, n31402, n31404, n31406, n31408, n31410, n31413, n31415,
         n31417, n31419, n31421, n31423, n31425, n31427, n31429, n31431,
         n31433, n31435, n31437, n31439, n31441, n31443, n31445, n31447,
         n31449, n31452, n31454, n31456, n31458, n31460, n31462, n31464,
         n31466, n31468, n31470, n31472, n31474, n31476, n31478, n31480,
         n31482, n31484, n31486, n31488, n31490, n31492, n31494, n31496,
         n31498, n31500, n31502, n31504, n31506, n31508, n31510, n31512,
         n31514, n31516, n31518, n31520, n31522, n31524, n31526, n31528,
         n31530, n31532, n31534, n31536, n31538, n31540, n31542, n31544,
         n31546, n31548, n31550, n31552, n31554, n31556, n31558, n31560,
         n31562, n31564, n31566, n31568, n31570, n31572, n31574, n31576,
         n31578, n31580, n31582, n31584, n31586, n31588, n31590, n31592,
         n31594, n31596, n31598, n31600, n31602, n31604, n31606, n31608,
         n31610, n31612, n31614, n31616, n31618, n31620, n31622, n31624,
         n31626, n31628, n31630, n31632, n31634, n31636, n31638, n31640,
         n31642, n31644, n31646, n31648, n31650, n31652, n31654, n31656,
         n31658, n31660, n31662, n31664, n31666, n31668, n31670, n31672,
         n31674, n31676, n31678, n31680, n31682, n31684, n31686, n31688,
         n31690, n31692, n31694, n31696, n31698, n31700, n31702, n31704,
         n31706, n31708, n31710, n31712, n31714, n31716, n31718, n31720,
         n31722, n31724, n31726, n31728, n31730, n31732, n31734, n31736,
         n31738, n31740, n31742, n31745, n31747, n31749, n31751, n31753,
         n31755, n31757, n31759, n31761, n31763, n31765, n31767, n31769,
         n31771, n31773, n31775, n31777, n31779, n31781, n31783, n31785,
         n31787, n31789, n31791, n31793, n31795, n31797, n31799, n31801,
         n31803, n31805, n31807, n31809, n31811, n31813, n31815, n31817,
         n31819, n31821, n31823, n31825, n31827, n31829, n31831, n31833,
         n31835, n31837, n31839, n31841, n31843, n31845, n31847, n31849,
         n31851, n31853, n31855, n31857, n31859, n31861, n31863, n31865,
         n31867, n31869, n31871, n31873, n31875, n31877, n31879, n31881,
         n31883, n31885, n31887, n31889, n31891, n31893, n31895, n31897,
         n31899, n31901, n31903, n31905, n31907, n31909, n31911, n31913,
         n31915, n31917, n31919, n31921, n31923, n31925, n31927, n31929,
         n31931, n31933, n31935, n31937, n31939, n31941, n31943, n31945,
         n31947, n31949, n31951, n31953, n31955, n31957, n31959, n31961,
         n31963, n31965, n31967, n31969, n31971, n31973, n31975, n31977,
         n31979, n31981, n31983, n31985, n31987, n31989, n31991, n31993,
         n31995, n31997, n31999, n32002, n32004, n32006, n32008, n32010,
         n32012, n32014, n32016, n32018, n32020, n32022, n32024, n32026,
         n32028, n32030, n32032, n32034, n32036, n32038, n32040, n32042,
         n32044, n32046, n32048, n32050, n32052, n32054, n32056, n32058,
         n32060, n32062, n32064, n32066, n32068, n32070, n32072, n32074,
         n32076, n32078, n32080, n32082, n32084, n32086, n32088, n32090,
         n32092, n32094, n32096, n32098, n32100, n32102, n32104, n32106,
         n32108, n32110, n32112, n32114, n32116, n32118, n32120, n32122,
         n32124, n32126, n32128, n32130, n32132, n32134, n32136, n32138,
         n32140, n32142, n32144, n32146, n32148, n32150, n32152, n32154,
         n32156, n32158, n32160, n32162, n32164, n32166, n32168, n32170,
         n32172, n32174, n32176, n32178, n32180, n32182, n32184, n32186,
         n32188, n32190, n32192, n32194, n32196, n32198, n32200, n32202,
         n32204, n32206, n32208, n32210, n32212, n32214, n32216, n32218,
         n32220, n32222, n32224, n32226, n32228, n32230, n32232, n32234,
         n32236, n32238, n32240, n32242, n32244, n32246, n32248, n32250,
         n32252, n32254, n32256, n32258, n32260, n32262, n32264, n32266,
         n32268, n32270, n32272, n32274, n32276, n32278, n32280, n32282,
         n32284, n32286, n32288, n32290, n32292, n32294, n32296, n32298,
         n32300, n32302, n32304, n32306, n32308, n32310, n32312, n32314,
         n32316, n32318, n32320, n32322, n32324, n32326, n32328, n32330,
         n32332, n32334, n32336, n32338, n32340, n32342, n32344, n32346,
         n32348, n32350, n32352, n32354, n32356, n32358, n32360, n32362,
         n32364, n32366, n32368, n32370, n32372, n32374, n32376, n32378,
         n32380, n32382, n32384, n32386, n32388, n32390, n32392, n32394,
         n32396, n32398, n32400, n32402, n32404, n32406, n32408, n32410,
         n32412, n32414, n32416, n32418, n32420, n32422, n32424, n32426,
         n32428, n32430, n32432, n32434, n32436, n32438, n32440, n32442,
         n32444, n32446, n32448, n32450, n32452, n32454, n32456, n32458,
         n32460, n32462, n32464, n32466, n32468, n32470, n32472, n32474,
         n32476, n32478, n32480, n32482, n32484, n32486, n32488, n32490,
         n32492, n32494, n32496, n32498, n32500, n32502, n32504, n32506,
         n32508, n32510, n32512, n32514, n32516, n32518, n32520, n32522,
         n32524, n32526, n32528, n32530, n32532, n32534, n32536, n32538,
         n32540, n32542, n32544, n32546, n32548, n32550, n32552, n32554,
         n32556, n32558, n32560, n32562, n32564, n32566, n32568, n32570,
         n32572, n32574, n32576, n32578, n32580, n32582, n32584, n32586,
         n32588, n32590, n32592, n32594, n32596, n32598, n32600, n32602,
         n32604, n32606, n32608, n32610, n32612, n32614, n32616, n32618,
         n32620, n32622, n32624, n32626, n32628, n32630, n32632, n32634,
         n32636, n32638, n32640, n32642, n32644, n32646, n32648, n32650,
         n32652, n32654, n32656, n32658, n32660, n32662, n32664, n32666,
         n32668, n32670, n32672, n32674, n32676, n32678, n32680, n32682,
         n32684, n32686, n32688, n32690, n32692, n32694, n32696, n32698,
         n32700, n32702, n32704, n32706, n32708, n32710, n32712, n32714,
         n32716, n32718, n32720, n32722, n32724, n32726, n32728, n32730,
         n32732, n32734, n32736, n32738, n32740, n32742, n32744, n32746,
         n32748, n32750, n32752, n32754, n32756, n32758, n32760, n32762,
         n32764, n32766, n32768, n32770, n32772, n32774, n32776, n32778,
         n32780, n32782, n32784, n32786, n32788, n32790, n32792, n32794,
         n32796, n32798, n32800, n32802, n32804, n32806, n32808, n32810,
         n32812, n32814, n32816, n32818, n32821, n32823, n32825, n32827,
         n32829, n32831, n32833, n32835, n32837, n32839, n32841, n32843,
         n32845, n32847, n32849, n32851, n32853, n32855, n32857, n32859,
         n32861, n32863, n32865, n32867, n32869, n32871, n32873, n32875,
         n32877, n32879, n32881, n32883, n32885, n32887, n32889, n32891,
         n32893, n32895, n32897, n32899, n32901, n32903, n32905, n32907,
         n32909, n32911, n32913, n32915, n32917, n32919, n32921, n32923,
         n32925, n32927, n32929, n32931, n32933, n32935, n32937, n32939,
         n32941, n32943, n32945, n32947, n32949, n32951, n32953, n32955,
         n32957, n32959, n32961, n32963, n32965, n32967, n32969, n32971,
         n32973, n32975, n32977, n32979, n32981, n32983, n32985, n32987,
         n32989, n32991, n32993, n32995, n32997, n32999, n33001, n33003,
         n33005, n33007, n33009, n33011, n33013, n33015, n33017, n33019,
         n33021, n33023, n33025, n33027, n33029, n33031, n33033, n33035,
         n33037, n33039, n33041, n33043, n33045, n33047, n33049, n33051,
         n33053, n33055, n33057, n33059, n33061, n33063, n33065, n33067,
         n33069, n33071, n33073, n33075, n33077, n33079, n33081, n33083,
         n33085, n33087, n33089, n33091, n33093, n33095, n33097, n33099,
         n33101, n33103, n33105, n33107, n33109, n33111, n33113, n33115,
         n33117, n33119, n33121, n33123, n33125, n33127, n33129, n33131,
         n33133, n33135, n33137, n33139, n33141, n33143, n33145, n33147,
         n33149, n33151, n33153, n33155, n33157, n33159, n33161, n33163,
         n33165, n33167, n33169, n33171, n33173, n33175, n33177, n33179,
         n33181, n33183, n33185, n33187, n33189, n33191, n33193, n33195,
         n33197, n33199, n33201, n33203, n33205, n33207, n33209, n33211,
         n33213, n33215, n33217, n33219, n33221, n33223, n33225, n33227,
         n33229, n33231, n33233, n33235, n33237, n33239, n33241, n33243,
         n33245, n33247, n33249, n33251, n33253, n33255, n33257, n33259,
         n33261, n33263, n33265, n33267, n33269, n33271, n33273, n33275,
         n33277, n33279, n33281, n33283, n33285, n33287, n33289, n33291,
         n33293, n33295, n33297, n33299, n33301, n33303, n33305, n33307,
         n33309, n33311, n33313, n33315, n33317, n33319, n33321, n33323,
         n33325, n33327, n33329, n33331, n33333, n33335, n33337, n33339,
         n33341, n33343, n33345, n33347, n33349, n33351, n33353, n33355,
         n33357, n33359, n33361, n33363, n33365, n33367, n33369, n33371,
         n33373, n33375, n33377, n33379, n33381, n33383, n33385, n33387,
         n33389, n33391, n33393, n33395, n33397, n33399, n33401, n33403,
         n33405, n33407, n33409, n33411, n33413, n33415, n33417, n33419,
         n33421, n33423, n33425, n33427, n33429, n33431, n33433, n33435,
         n33437, n33439, n33441, n33443, n33445, n33447, n33449, n33451,
         n33453, n33455, n33457, n33459, n33461, n33463, n33465, n33467,
         n33469, n33471, n33473, n33475, n33477, n33479, n33481, n33483,
         n33485, n33487, n33489, n33491, n33493, n33495, n33497, n33499,
         n33501, n33503, n33505, n33507, n33509, n33511, n33513, n33515,
         n33517, n33519, n33521, n33523, n33525, n33527, n33529, n33531,
         n33533, n33535, n33537, n33539, n33541, n33543, n33545, n33547,
         n33549, n33551, n33553, n33555, n33557, n33559, n33561, n33563,
         n33565, n33567, n33569, n33571, n33573, n33575, n33577, n33579,
         n33581, n33583, n33585, n33587, n33589, n33591, n33593, n33595,
         n33597, n33599, n33601, n33603, n33605, n33607, n33609, n33611,
         n33613, n33615, n33617, n33619, n33621, n33623, n33625, n33627,
         n33629, n33631, n33633, n33635, n33637, n33639, n33641, n33643,
         n33645, n33647, n33649, n33651, n33653, n33655, n33657, n33659,
         n33661, n33663, n33665, n33667, n33669, n33671, n33673, n33675,
         n33677, n33679, n33681, n33683, n33685, n33687, n33689, n33691,
         n33693, n33695, n33697, n33699, n33701, n33703, n33705, n33707,
         n33709, n33711, n33713, n33715, n33717, n33719, n33721, n33723,
         n33725, n33727, n33729, n33731, n33733, n33735, n33737, n33739,
         n33741, n33743, n33745, n33747, n33749, n33751, n33753, n33755,
         n33757, n33759, n33761, n33763, n33765, n33767, n33769, n33771,
         n33773, n33775, n33777, n33779, n33781, n33783, n33785, n33787,
         n33789, n33791, n33793, n33795, n33797, n33799, n33801, n33803,
         n33805, n33807, n33809, n33811, n33813, n33815, n33817, n33819,
         n33821, n33823, n33825, n33827, n33829, n33831, n33833, n33835,
         n33837, n33839, n33841, n33843, n33845, n33847, n33849, n33851,
         n33853, n33855, n33857, n33859, n33861, n33863, n33865, n33867,
         n33869, n33871, n33873, n33875, n33877, n33879, n33881, n33883,
         n33885, n33887, n33889, n33891, n33893, n33895, n33897, n33899,
         n33901, n33903, n33905, n33907, n33909, n33911, n33913, n33915,
         n33917, n33919, n56492, n56498, n56495, n56496, n56494, n56382,
         n33936, n33938, n33941, n33943, n64221, n64222, n64223, n64224,
         n64225, n64226, n64227, n64228, n64229, n64230, n64231, n64232,
         n64233, n64234, n64235, n64236, n64237, n64238, n64239, n64240,
         n64241, n64242, n64243, n64244, n64245, n64246, n64247, n64248,
         n64249, n64250, n64251, n64252, n64253, n64254, n64255, n64256,
         n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264,
         n64265, n64266, n64267, n64268, n64269, n64270, n64271, n64272,
         n64273, n64274, n64275, n64276, n64277, n64278, n64279, n64280,
         n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288,
         n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296,
         n64297, n64298, n64299, n64300, n64301, n64302, n64303, n64304,
         n64305, n64306, n64307, n64308, n64309, n64310, n64311, n64312,
         n64313, n64314, n64315, n64316, n64317, n64318, n64319, n64320,
         n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328,
         n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336,
         n64337, n64338, n64339, n64340, n64341, n64342, n64343, n64344,
         n64345, n64346, n64347, n64348, n64349, n64350, n64351, n64352,
         n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360,
         n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368,
         n64369, n64370, n64371, n64372, n64373, n64374, n64375, n64376,
         n64377, n64378, n64379, n64380, n64381, n64382, n64383, n64384,
         n64385, n64386, n64387, n64388, n64389, n64390, n64391, n64392,
         n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400,
         n64401, n64402, n64403, n64404, n64405, n64406, n64407, n64408,
         n64409, n64410, n64411, n64412, n64413, n64414, n64415, n64416,
         n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424,
         n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432,
         n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440,
         n64441, n64442, n64443, n64444, n64445, n64446, n64447, n64448,
         n64449, n64450, n64451, n64452, n64453, n64454, n64455, n64456,
         n64457, n64458, n64459, n64460, n64462, n64463, n64465, n64466,
         n64467, n34470, n34472, n34474, n34476, n34478, n34480, n34482,
         n34484, n34486, n34488, n34490, n34492, n34494, n34496, n34498,
         n34500, n34502, n34504, n34506, n34508, n34510, n34512, n34514,
         n34516, n34518, n34520, n34522, n34524, n34526, n34528, n34530,
         n34532, n34534, n34536, n34538, n34540, n34542, n34544, n34546,
         n34548, n34550, n34552, n34554, n34556, n34558, n34560, n34562,
         n34564, n34566, n34568, n34570, n34572, n34574, n34576, n34578,
         n34580, n34582, n34584, n34586, n34588, n34590, n34592, n34594,
         n34596, n34598, n34600, n34602, n34604, n34606, n34608, n34610,
         n34612, n34614, n34616, n34618, n34620, n34622, n34624, n34626,
         n34628, n34630, n34632, n34634, n34636, n34638, n34640, n34642,
         n34644, n34646, n34648, n34650, n34652, n34654, n34656, n34658,
         n34660, n34662, n34664, n34666, n34668, n34670, n34672, n34674,
         n34676, n34678, n34680, n34682, n34684, n34686, n34688, n34690,
         n34692, n34694, n34696, n34698, n34700, n34702, n34704, n34706,
         n34708, n34710, n34712, n34714, n34716, n34718, n34720, n34722,
         n34724, n34726, n34728, n34730, n34732, n34734, n34736, n34738,
         n34740, n34742, n34744, n34746, n34748, n34750, n34752, n34754,
         n34756, n34758, n34760, n34762, n34764, n34766, n34768, n34770,
         n34772, n34774, n34776, n34778, n34780, n34782, n34784, n34786,
         n34788, n34790, n34792, n34794, n34796, n34798, n34800, n34802,
         n34804, n34806, n34808, n34810, n34812, n34814, n34816, n34818,
         n34820, n34822, n34824, n34826, n34828, n34830, n34832, n34834,
         n34836, n34838, n34840, n34842, n34844, n34846, n34848, n34850,
         n34852, n34854, n34856, n34858, n34860, n34862, n34864, n34866,
         n34868, n34870, n34872, n34874, n34876, n34878, n34880, n34882,
         n34884, n34886, n34888, n34890, n34892, n34894, n34896, n34898,
         n34900, n34902, n34904, n34906, n34908, n34910, n34912, n34914,
         n34916, n34918, n34920, n34922, n34924, n34926, n34928, n34930,
         n34932, n34934, n34936, n34938, n34940, n34942, n34944, n34946,
         n34948, n34950, n34952, n34954, n34956, n34958, n34960, n34962,
         n34964, n34966, n34968, n34970, n34972, n34974, n34976, n34978,
         n34980, n34982, n34984, n34986, n34988, n34990, n34992, n34994,
         n34996, n34998, n35000, n35002, n35004, n35006, n35008, n35010,
         n35012, n35014, n35016, n35018, n35020, n35022, n35024, n35026,
         n35028, n35030, n35032, n35034, n35036, n35038, n35040, n35042,
         n35044, n35046, n35048, n35050, n35052, n35054, n35056, n35058,
         n35060, n35062, n35064, n35066, n35068, n35070, n35072, n35074,
         n35076, n35078, n35080, n35082, n35084, n35086, n35088, n35090,
         n35092, n35094, n35096, n35098, n35100, n35102, n35104, n35106,
         n35108, n35110, n35112, n35114, n35116, n35118, n35120, n35122,
         n35124, n35126, n35128, n35130, n35132, n35134, n35136, n35138,
         n35140, n35142, n35144, n35146, n35148, n35150, n35152, n35154,
         n35156, n35158, n35160, n35162, n35164, n35166, n35168, n35170,
         n35172, n35174, n35176, n35178, n35180, n35182, n35184, n35186,
         n35188, n35190, n35192, n35194, n35196, n35198, n35200, n35202,
         n35204, n35206, n35208, n35210, n35212, n35214, n35216, n35218,
         n35220, n35222, n35224, n35226, n35228, n35230, n35232, n35234,
         n35236, n35238, n35240, n35242, n35244, n35246, n35248, n35250,
         n35252, n35254, n35256, n35258, n35260, n35262, n35264, n35266,
         n35268, n35270, n35272, n35274, n35276, n35278, n35280, n35282,
         n35284, n35286, n35288, n35290, n35292, n35294, n35296, n35298,
         n35300, n35302, n35304, n35306, n35308, n35310, n35312, n35314,
         n35316, n35318, n35320, n35322, n35324, n35326, n35328, n35330,
         n35332, n35334, n35336, n35338, n35340, n35342, n35344, n35346,
         n35348, n35350, n35352, n35354, n35356, n35358, n35360, n35362,
         n35364, n35366, n35368, n35370, n35372, n35374, n35376, n35378,
         n35380, n35382, n35384, n35386, n35388, n35390, n35392, n35394,
         n35396, n35398, n35400, n35402, n35404, n35406, n35408, n35410,
         n35412, n35414, n35416, n35418, n35420, n35422, n35424, n35426,
         n35428, n35430, n35432, n35434, n35436, n35438, n35440, n35442,
         n35444, n35446, n35448, n35450, n35452, n35454, n35456, n35458,
         n35460, n35462, n35464, n35466, n35468, n35470, n35472, n35474,
         n35476, n35478, n35480, n35482, n35484, n35486, n35488, n35490,
         n35492, n35494, n35496, n35498, n35500, n35502, n35504, n35506,
         n35508, n35510, n35512, n35514, n35516, n35518, n35520, n35522,
         n35524, n35526, n35528, n35530, n35532, n35534, n35536, n35538,
         n35540, n35542, n35544, n35546, n35548, n35550, n35552, n35554,
         n35556, n35558, n35560, n35562, n35564, n35566, n35568, n35570,
         n35572, n35574, n35576, n35578, n35580, n35582, n35584, n35586,
         n35588, n35590, n35592, n35594, n35596, n35598, n35600, n35602,
         n35604, n35606, n35608, n35610, n35612, n35614, n35616, n35618,
         n35620, n35622, n35624, n35626, n35628, n35630, n35632, n35634,
         n35636, n35638, n35640, n35642, n35644, n35646, n35648, n35650,
         n35652, n35654, n35656, n35658, n35660, n35662, n35664, n35666,
         n35668, n35670, n35672, n35674, n35676, n35678, n35680, n35682,
         n35684, n35686, n35688, n35690, n35692, n35694, n35696, n35698,
         n35700, n35702, n35704, n35706, n35708, n35710, n35712, n35714,
         n35716, n35718, n35720, n35722, n35724, n35726, n35728, n35730,
         n35732, n35734, n35736, n35738, n35740, n35742, n35744, n35746,
         n35748, n35750, n35752, n35754, n35756, n35758, n35760, n35762,
         n35764, n35766, n35768, n35770, n35772, n35774, n35776, n35778,
         n35780, n35782, n35784, n35786, n35788, n35790, n35792, n35794,
         n35796, n35798, n35800, n35802, n35804, n35806, n35808, n35810,
         n35812, n35814, n35816, n35818, n35820, n35822, n35824, n35826,
         n35828, n35830, n35832, n35834, n35836, n35838, n35840, n35842,
         n35844, n35846, n35848, n35850, n35852, n35854, n35856, n35858,
         n35860, n35862, n35864, n35866, n35868, n35870, n35872, n35874,
         n35876, n64213, n64214, n64210, n64208, n64209, n64205, n64206,
         n64207, n64201, n64202, n64203, n64204, n64197, n64198, n64199,
         n64200, n64193, n64194, n64195, n64196, n64189, n64190, n64191,
         n64192, n64185, n64186, n64187, n64188, n64181, n64182, n64183,
         n64184, n64177, n64178, n64179, n64180, n64173, n64174, n64175,
         n64176, n64169, n64170, n64171, n64172, n64165, n64166, n64167,
         n64168, n64161, n64162, n64163, n64164, n64157, n64158, n64159,
         n64160, n64153, n64154, n64155, n64156, n64149, n64150, n64151,
         n64152, n64145, n64146, n64147, n64148, n64141, n64142, n64143,
         n64144, n64137, n64138, n64139, n64140, n64133, n64134, n64135,
         n64136, n64129, n64130, n64131, n64132, n64125, n64126, n64127,
         n64128, n36059, n36061, n36063, n36065, n36067, n36069, n36071,
         n36073, n36075, n36077, n36079, n36081, n36083, n36085, n36087,
         n36089, n36091, n36093, n36095, n36097, n36099, n36101, n36103,
         n36105, n36107, n36109, n36111, n36113, n36115, n36117, n36119,
         n36121, n36123, n36125, n36127, n36129, n36131, n36133, n36135,
         n36137, n36139, n36141, n36143, n36145, n36147, n36149, n36151,
         n36153, n36155, n36157, n36159, n36161, n36163, n36165, n36167,
         n36169, n36171, n36173, n36175, n36177, n36179, n36181, n36183,
         n36185, n36187, n36189, n36191, n36193, n36195, n36197, n36199,
         n36201, n36203, n36205, n36207, n36209, n36211, n36213, n36215,
         n36217, n36219, n36221, n36223, n36225, n36227, n36229, n36231,
         n36233, n36235, n36237, n36239, n36241, n36243, n36245, n36247,
         n36249, n36251, n36253, n36255, n36257, n36259, n36261, n36263,
         n36265, n36267, n36269, n36271, n36273, n36275, n36277, n36279,
         n36281, n36283, n36285, n36287, n36289, n36291, n36293, n36295,
         n36297, n36299, n36301, n36303, n36305, n36307, n36309, n36311,
         n36313, n36315, n36317, n36319, n36321, n36323, n36325, n36327,
         n36329, n36331, n36333, n36335, n36337, n36339, n36341, n36343,
         n36345, n36347, n36349, n36351, n36353, n36355, n36357, n36359,
         n36361, n36363, n36365, n36367, n36369, n36371, n36373, n36375,
         n36377, n36379, n36381, n36383, n36385, n36387, n36389, n36391,
         n36393, n36395, n36397, n36399, n36401, n36403, n36405, n36407,
         n36409, n36411, n36413, n36415, n36417, n36419, n36421, n36423,
         n36425, n36427, n36429, n36431, n36433, n36435, n36437, n36439,
         n36441, n36443, n36445, n36447, n36449, n36451, n36453, n36455,
         n36457, n36459, n36461, n36463, n36465, n36467, n36469, n36471,
         n36473, n36475, n36477, n36479, n36481, n36483, n36485, n36487,
         n36489, n36491, n36493, n36495, n36497, n36499, n36501, n36503,
         n36505, n36507, n36509, n36511, n36513, n36515, n36517, n36519,
         n36521, n36523, n36525, n36527, n36529, n36531, n36533, n36535,
         n36537, n36539, n36541, n36543, n36545, n36547, n36549, n36551,
         n36553, n36555, n36557, n36559, n36561, n36563, n36565, n36567,
         n36569, n36571, n36573, n36575, n36577, n36579, n36581, n36583,
         n36585, n36587, n36589, n36591, n36593, n36595, n36597, n36599,
         n36601, n36603, n36605, n36607, n36609, n36611, n36613, n36615,
         n36617, n36619, n36621, n36623, n36625, n36627, n36629, n36631,
         n36633, n36635, n36637, n36639, n36641, n36643, n36645, n36647,
         n36649, n36651, n36653, n36655, n36657, n36659, n36661, n36663,
         n36665, n36667, n36669, n36671, n36673, n36675, n36677, n36679,
         n36681, n36683, n36685, n36687, n36689, n36691, n36693, n36695,
         n36697, n36699, n36701, n36703, n36705, n36707, n36709, n36711,
         n36713, n36715, n36717, n36719, n36721, n36723, n36725, n36727,
         n36729, n36731, n36733, n36735, n36737, n36739, n36741, n36743,
         n36745, n36747, n36749, n36751, n36753, n36755, n36757, n36759,
         n36761, n36763, n36765, n36767, n36769, n36771, n36773, n36775,
         n36777, n36779, n36781, n36783, n36785, n36787, n36789, n36791,
         n36793, n36795, n36797, n36799, n36801, n36803, n36805, n36807,
         n36809, n36811, n36813, n36815, n36817, n36819, n36821, n36823,
         n36825, n36827, n36829, n36831, n36833, n36835, n36837, n36839,
         n36841, n36843, n36845, n36847, n36849, n36851, n36853, n36855,
         n36857, n36859, n36861, n36863, n36865, n36867, n36869, n36871,
         n36873, n36875, n36877, n36879, n36881, n36883, n36885, n36887,
         n36889, n36891, n36893, n36895, n36897, n36899, n36901, n36903,
         n36905, n36907, n36909, n36911, n36913, n36915, n36917, n36919,
         n36921, n36923, n36925, n36927, n36929, n36931, n36933, n36935,
         n36937, n36939, n36941, n36943, n36945, n36947, n36949, n36951,
         n36953, n36955, n36957, n36959, n36961, n36963, n36965, n36967,
         n36969, n36971, n36973, n36975, n36977, n36979, n36981, n36983,
         n36985, n36987, n36989, n36991, n36993, n36995, n36997, n36999,
         n37001, n37003, n37005, n37007, n37009, n37011, n37013, n37015,
         n37017, n37019, n37021, n37023, n37025, n37027, n37029, n37031,
         n37033, n37035, n37037, n37039, n37041, n37043, n37045, n37047,
         n37049, n37051, n37053, n37055, n37057, n37059, n37061, n37063,
         n37065, n37067, n37069, n37071, n37073, n37075, n37077, n37079,
         n37081, n37083, n37085, n37087, n37089, n37091, n37093, n37095,
         n37097, n37099, n37101, n37103, n37105, n37107, n37109, n37111,
         n37113, n37115, n37117, n37119, n37121, n37123, n37125, n37127,
         n37129, n37131, n37133, n37135, n37137, n37139, n37141, n37143,
         n37145, n37147, n37149, n37151, n37153, n37155, n37157, n37159,
         n37161, n37163, n37165, n37167, n37169, n37171, n37173, n37175,
         n37177, n37179, n37181, n37183, n37185, n37187, n37189, n37191,
         n37193, n37195, n37197, n37199, n37201, n37203, n37205, n37207,
         n37209, n37211, n37213, n37215, n37217, n37219, n37221, n37223,
         n37225, n37227, n37229, n37231, n37233, n37235, n37237, n37239,
         n37241, n37243, n37245, n37247, n37249, n37251, n37253, n37255,
         n37257, n37259, n37261, n37263, n37265, n37267, n37269, n37271,
         n37273, n37275, n37277, n37279, n37281, n37283, n37285, n37287,
         n37289, n37291, n37293, n37295, n37297, n37299, n37301, n37303,
         n37305, n37307, n37309, n37311, n37313, n37315, n37317, n37319,
         n37321, n37323, n37325, n37327, n37329, n37331, n37333, n37335,
         n37337, n37339, n37341, n37343, n37345, n37347, n37349, n37351,
         n37353, n37355, n37357, n37359, n37361, n37363, n37365, n37367,
         n37369, n37371, n37373, n37375, n37377, n37379, n37381, n37383,
         n37385, n37387, n37389, n37391, n37393, n37395, n37397, n37399,
         n37401, n37403, n37405, n37407, n37409, n37411, n37413, n37415,
         n37417, n37419, n37421, n37423, n37425, n37427, n37429, n37431,
         n37433, n37435, n37437, n37439, n37441, n37443, n37445, n37447,
         n37449, n37451, n37453, n37455, n37457, n37459, n37461, n37463,
         n37465, n37467, n37469, n37471, n37473, n37475, n37477, n37479,
         n37481, n37483, n37485, n37487, n37489, n37491, n37493, n37495,
         n37497, n37499, n37501, n37503, n37505, n37507, n37509, n37511,
         n37513, n37515, n37517, n37519, n37521, n37523, n37525, n37527,
         n37529, n37531, n37533, n37535, n37537, n37539, n37541, n37543,
         n37545, n37547, n37549, n37551, n37553, n37555, n37557, n37559,
         n37561, n37563, n37565, n37567, n37569, n37571, n37573, n37575,
         n37577, n37579, n37581, n37583, n37585, n37587, n37589, n37591,
         n37593, n37595, n37597, n37599, n37601, n37603, n37605, n37607,
         n37609, n37611, n37613, n37615, n37617, n37619, n37621, n37623,
         n37625, n37627, n37629, n37631, n37633, n37635, n37637, n37639,
         n37641, n37643, n37645, n37647, n37649, n37651, n37653, n37655,
         n37657, n37659, n37661, n37663, n37665, n37667, n37669, n37671,
         n37673, n37675, n37677, n37679, n37681, n37683, n37685, n37687,
         n37689, n37691, n37693, n37695, n37697, n37699, n37701, n37703,
         n37705, n37707, n37709, n37711, n37713, n37715, n37717, n37719,
         n37721, n37723, n37725, n37727, n37729, n37731, n37733, n37735,
         n37737, n37739, n37741, n37743, n37745, n37747, n37749, n37751,
         n37753, n37755, n37757, n37759, n37761, n37763, n37765, n37767,
         n37769, n37771, n37773, n37775, n37777, n37779, n37781, n37783,
         n37785, n37787, n37789, n37791, n37793, n37795, n37797, n37799,
         n37801, n37803, n37805, n37807, n37809, n37811, n37813, n37815,
         n37817, n37819, n37821, n37823, n37825, n37827, n37829, n37831,
         n37833, n37835, n37837, n37839, n37841, n37843, n37845, n37847,
         n37849, n37851, n37853, n37855, n37857, n37859, n37861, n37863,
         n37865, n37867, n37869, n37871, n37873, n37875, n37877, n37879,
         n37881, n37883, n37885, n37887, n37889, n37891, n37893, n37895,
         n37897, n37899, n37901, n37903, n37905, n37907, n37909, n37911,
         n37913, n37915, n37917, n37919, n37921, n37923, n37925, n37927,
         n37929, n37931, n37933, n37935, n37937, n37939, n37941, n37943,
         n37945, n37947, n37949, n37951, n37953, n37955, n37957, n37959,
         n37961, n37963, n37965, n37967, n37969, n37971, n37973, n37975,
         n37977, n37979, n37981, n37983, n37985, n37987, n37989, n37991,
         n37993, n37995, n37997, n37999, n38001, n38003, n38005, n38007,
         n38009, n38011, n38013, n38015, n38017, n38019, n38021, n38023,
         n38025, n38027, n38029, n38031, n38033, n38035, n38037, n38039,
         n38041, n38043, n38045, n38047, n38049, n38051, n38053, n38055,
         n38057, n38059, n38061, n38063, n38065, n38067, n38069, n38071,
         n38073, n38075, n38077, n38079, n38081, n38083, n38085, n38087,
         n38089, n38091, n38093, n38095, n38097, n38099, n38101, n38103,
         n38105, n38107, n38109, n38111, n38113, n38115, n38117, n38119,
         n38121, n38123, n38125, n38127, n38129, n38131, n38133, n38135,
         n38137, n38139, n38141, n38143, n38145, n38147, n38149, n38151,
         n38153, n38155, n38157, n38159, n38161, n38163, n38165, n38167,
         n38169, n38171, n38173, n38175, n38177, n38179, n38181, n38183,
         n38185, n38187, n38189, n38191, n38193, n38195, n38197, n38199,
         n38201, n38203, n38205, n38207, n38209, n38211, n38213, n38215,
         n38217, n38219, n38221, n38223, n38225, n38227, n38229, n38231,
         n38233, n38235, n38237, n38239, n38241, n38243, n38245, n38247,
         n38249, n38251, n38253, n38255, n38257, n38259, n38261, n38263,
         n38265, n38267, n38269, n38271, n38273, n38275, n38277, n38279,
         n38281, n38283, n38285, n38287, n38289, n38291, n38293, n38295,
         n38297, n38299, n38301, n38303, n38305, n38307, n38309, n38311,
         n38313, n38315, n38317, n38319, n38321, n38323, n38325, n38327,
         n38329, n38331, n38333, n38335, n38337, n38339, n38341, n38343,
         n38345, n38347, n38349, n38351, n38353, n38355, n38357, n38359,
         n38361, n38363, n38365, n38367, n38369, n38371, n38373, n38375,
         n38377, n38379, n38381, n38383, n38385, n38387, n38389, n38391,
         n38393, n38395, n38397, n38399, n38401, n38403, n38405, n38407,
         n38409, n38411, n38413, n38415, n38417, n38419, n38421, n38423,
         n38425, n38427, n38429, n38431, n38433, n38435, n38437, n38439,
         n38441, n38443, n38445, n38447, n38449, n38451, n38453, n38455,
         n38457, n38459, n38461, n38463, n38465, n38467, n38469, n38471,
         n38473, n38475, n38477, n38479, n38481, n38483, n38485, n38487,
         n38489, n38491, n38493, n38495, n38497, n38499, n38501, n38503,
         n38505, n38507, n38509, n38511, n38513, n38515, n38517, n38519,
         n38521, n38523, n38525, n38527, n38529, n38531, n38533, n38535,
         n38537, n38539, n38541, n38543, n38545, n38547, n38549, n38551,
         n38553, n38555, n38557, n38559, n38561, n38563, n38565, n38567,
         n38569, n38571, n38573, n38575, n38577, n38579, n38581, n38583,
         n38585, n38587, n38589, n38591, n38593, n38595, n38597, n38599,
         n38601, n38603, n38605, n38607, n38609, n38611, n38613, n38615,
         n38617, n38619, n38621, n38623, n38625, n38627, n38629, n38631,
         n38633, n38635, n38637, n38639, n38641, n38643, n38645, n38647,
         n38649, n38651, n38653, n38655, n38657, n38659, n38661, n38663,
         n38665, n38667, n38669, n38671, n38673, n38675, n38677, n38679,
         n38681, n38683, n38685, n38687, n38689, n38691, n38693, n38695,
         n38697, n38699, n38701, n38703, n38705, n38707, n38709, n38711,
         n38713, n38715, n38717, n38719, n38721, n38723, n38725, n38727,
         n38729, n38731, n38733, n38735, n38737, n38739, n38741, n38743,
         n38745, n38747, n38749, n38751, n38753, n38755, n38757, n38759,
         n38761, n38763, n38765, n38767, n38769, n38771, n38773, n38775,
         n38777, n38779, n38781, n38783, n38785, n38787, n38789, n38791,
         n38793, n38795, n38797, n38799, n38801, n38803, n38805, n38807,
         n38809, n38811, n38813, n38815, n38817, n38819, n38821, n38823,
         n38825, n38827, n38829, n38831, n38833, n38835, n38837, n38839,
         n38841, n38843, n38845, n38847, n38849, n38851, n38853, n38855,
         n38857, n38859, n38861, n38863, n38865, n38867, n38869, n38871,
         n38873, n38875, n38877, n38879, n38881, n38883, n38885, n38887,
         n38889, n38891, n38893, n38895, n38897, n38899, n38901, n38903,
         n38905, n38907, n38909, n38911, n38913, n38915, n38917, n38919,
         n38921, n38923, n38925, n38927, n38929, n38931, n38933, n38935,
         n38937, n38939, n38941, n38943, n38945, n38947, n38949, n38951,
         n38953, n38955, n38957, n38959, n38961, n38963, n38965, n38967,
         n38969, n38971, n38973, n38975, n38977, n38979, n38981, n38983,
         n38985, n38987, n38989, n38991, n38993, n38995, n38997, n38999,
         n39001, n39003, n39005, n39007, n39009, n39011, n39013, n39015,
         n39017, n39019, n39021, n39023, n39025, n39027, n39029, n39031,
         n39033, n39035, n39037, n39039, n39041, n39043, n39045, n39047,
         n39049, n39051, n39053, n39055, n39057, n39059, n39061, n39063,
         n39065, n39067, n39069, n39071, n39073, n39075, n39077, n39079,
         n39081, n39083, n39085, n39087, n39089, n39091, n39093, n39095,
         n39097, n39099, n39101, n39103, n39105, n39107, n39109, n39111,
         n39113, n39115, n39117, n39119, n39121, n39123, n39125, n39127,
         n39129, n39131, n39133, n39135, n39137, n39139, n39141, n39143,
         n39145, n39147, n39149, n39151, n39153, n39155, n39157, n39159,
         n39161, n39163, n39165, n39167, n39169, n39171, n39173, n39175,
         n39177, n39179, n39181, n39183, n39185, n39187, n39189, n39191,
         n39193, n39195, n39197, n39199, n39201, n39203, n39205, n39207,
         n39209, n39211, n39213, n39215, n39217, n39219, n39221, n39223,
         n39225, n39227, n39229, n39231, n39233, n39235, n39237, n39239,
         n39241, n39243, n39245, n39247, n39249, n39251, n39253, n39255,
         n39257, n39259, n39261, n39263, n39265, n39267, n39269, n39271,
         n39273, n39275, n39277, n39279, n39281, n39283, n39285, n39287,
         n39289, n39291, n39293, n39295, n39297, n39299, n39301, n39303,
         n39305, n39307, n39309, n39311, n39313, n39315, n39317, n39319,
         n39321, n39323, n39325, n39327, n39329, n39331, n39333, n39335,
         n39337, n39339, n39341, n39343, n39345, n39347, n39349, n39351,
         n39353, n39355, n39357, n39359, n39361, n39363, n39365, n39367,
         n39369, n39371, n39373, n39375, n39377, n39379, n39381, n39383,
         n39385, n39387, n39389, n39391, n39393, n39395, n39397, n39399,
         n39401, n39403, n39405, n39407, n39409, n39411, n39413, n39415,
         n39417, n39419, n39421, n39423, n39425, n39427, n39429, n39431,
         n39433, n39435, n39437, n39439, n39441, n39443, n39445, n39447,
         n39449, n39451, n39453, n39455, n39457, n39459, n39461, n39463,
         n39465, n39467, n39469, n39471, n39473, n39475, n39477, n39479,
         n39481, n39483, n39485, n39487, n39489, n39491, n39493, n39495,
         n39497, n39499, n39501, n39503, n39505, n39515, n39522, n39524,
         n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533,
         n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541,
         n39542, n39543, n39544, n39545, n39546, n39547, n39548, n39549,
         n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557,
         n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565,
         n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573,
         n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581,
         n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589,
         n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597,
         n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605,
         n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613,
         n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621,
         n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629,
         n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637,
         n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645,
         n39646, n39647, n39648, n39649, n39653, n39655, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39694,
         n39696, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
         n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
         n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
         n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
         n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
         n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
         n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
         n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
         n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
         n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
         n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
         n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
         n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
         n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
         n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
         n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
         n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
         n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
         n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888,
         n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
         n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
         n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
         n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
         n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928,
         n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
         n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944,
         n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
         n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960,
         n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
         n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
         n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
         n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
         n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
         n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008,
         n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016,
         n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
         n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
         n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
         n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
         n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056,
         n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
         n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
         n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
         n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
         n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
         n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
         n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
         n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
         n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
         n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
         n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
         n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
         n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
         n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
         n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
         n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
         n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
         n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
         n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
         n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
         n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
         n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
         n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
         n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
         n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
         n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
         n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
         n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
         n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
         n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
         n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
         n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
         n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
         n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
         n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
         n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
         n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
         n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
         n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
         n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
         n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
         n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
         n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
         n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
         n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432,
         n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440,
         n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448,
         n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
         n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464,
         n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
         n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
         n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488,
         n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
         n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504,
         n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512,
         n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520,
         n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
         n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536,
         n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
         n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552,
         n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560,
         n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568,
         n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576,
         n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584,
         n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
         n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
         n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608,
         n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
         n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
         n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632,
         n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640,
         n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648,
         n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656,
         n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664,
         n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
         n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
         n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
         n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696,
         n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704,
         n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712,
         n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720,
         n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728,
         n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736,
         n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
         n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752,
         n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
         n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768,
         n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776,
         n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784,
         n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792,
         n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800,
         n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808,
         n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
         n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824,
         n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
         n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840,
         n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848,
         n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
         n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864,
         n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872,
         n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880,
         n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
         n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896,
         n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
         n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912,
         n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920,
         n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928,
         n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936,
         n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944,
         n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952,
         n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
         n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968,
         n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
         n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
         n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992,
         n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
         n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008,
         n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016,
         n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024,
         n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
         n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040,
         n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
         n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056,
         n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064,
         n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072,
         n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080,
         n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088,
         n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096,
         n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
         n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
         n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
         n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
         n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136,
         n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144,
         n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152,
         n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160,
         n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
         n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
         n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184,
         n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
         n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200,
         n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208,
         n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
         n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224,
         n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232,
         n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240,
         n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
         n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256,
         n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
         n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272,
         n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280,
         n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288,
         n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
         n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
         n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312,
         n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
         n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328,
         n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
         n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344,
         n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352,
         n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360,
         n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
         n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376,
         n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384,
         n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
         n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400,
         n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
         n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416,
         n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424,
         n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
         n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440,
         n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448,
         n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456,
         n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
         n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472,
         n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
         n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
         n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496,
         n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
         n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512,
         n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520,
         n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528,
         n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
         n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544,
         n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
         n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
         n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
         n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
         n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584,
         n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592,
         n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600,
         n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
         n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616,
         n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
         n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
         n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640,
         n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
         n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656,
         n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664,
         n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
         n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
         n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688,
         n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
         n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
         n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
         n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
         n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728,
         n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736,
         n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744,
         n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
         n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760,
         n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
         n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776,
         n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784,
         n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
         n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800,
         n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808,
         n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816,
         n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
         n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832,
         n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
         n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848,
         n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
         n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864,
         n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872,
         n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880,
         n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888,
         n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
         n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904,
         n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
         n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
         n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928,
         n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936,
         n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944,
         n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952,
         n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960,
         n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
         n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976,
         n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
         n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
         n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000,
         n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008,
         n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016,
         n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024,
         n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032,
         n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
         n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048,
         n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
         n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
         n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072,
         n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080,
         n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088,
         n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096,
         n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104,
         n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
         n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120,
         n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
         n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136,
         n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144,
         n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
         n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160,
         n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168,
         n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176,
         n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
         n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192,
         n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
         n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208,
         n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216,
         n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
         n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232,
         n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240,
         n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248,
         n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
         n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
         n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
         n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
         n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288,
         n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296,
         n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304,
         n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312,
         n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320,
         n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
         n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336,
         n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
         n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
         n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360,
         n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368,
         n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376,
         n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384,
         n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392,
         n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400,
         n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408,
         n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
         n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424,
         n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432,
         n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440,
         n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448,
         n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456,
         n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464,
         n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472,
         n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480,
         n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488,
         n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496,
         n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504,
         n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512,
         n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520,
         n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528,
         n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536,
         n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544,
         n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552,
         n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560,
         n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568,
         n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576,
         n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584,
         n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592,
         n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600,
         n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608,
         n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
         n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624,
         n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632,
         n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640,
         n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648,
         n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656,
         n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664,
         n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672,
         n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680,
         n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688,
         n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696,
         n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704,
         n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712,
         n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720,
         n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728,
         n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736,
         n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744,
         n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752,
         n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
         n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768,
         n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
         n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784,
         n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792,
         n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800,
         n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
         n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816,
         n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824,
         n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
         n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840,
         n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848,
         n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856,
         n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864,
         n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
         n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880,
         n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888,
         n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896,
         n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904,
         n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912,
         n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920,
         n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928,
         n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936,
         n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944,
         n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952,
         n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960,
         n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968,
         n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976,
         n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984,
         n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992,
         n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
         n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008,
         n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016,
         n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024,
         n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032,
         n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040,
         n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048,
         n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056,
         n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
         n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072,
         n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080,
         n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088,
         n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096,
         n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104,
         n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112,
         n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
         n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128,
         n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
         n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144,
         n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152,
         n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
         n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168,
         n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176,
         n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184,
         n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
         n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200,
         n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
         n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216,
         n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224,
         n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232,
         n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240,
         n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248,
         n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256,
         n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
         n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272,
         n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
         n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288,
         n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296,
         n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304,
         n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312,
         n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320,
         n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328,
         n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336,
         n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344,
         n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
         n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360,
         n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368,
         n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376,
         n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384,
         n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392,
         n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400,
         n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
         n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416,
         n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
         n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432,
         n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440,
         n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448,
         n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456,
         n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464,
         n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472,
         n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
         n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488,
         n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
         n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504,
         n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512,
         n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520,
         n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528,
         n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536,
         n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544,
         n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
         n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560,
         n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568,
         n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576,
         n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584,
         n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592,
         n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600,
         n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608,
         n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616,
         n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
         n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632,
         n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640,
         n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648,
         n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656,
         n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664,
         n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672,
         n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680,
         n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688,
         n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
         n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704,
         n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712,
         n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720,
         n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728,
         n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736,
         n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744,
         n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752,
         n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760,
         n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
         n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776,
         n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
         n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792,
         n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800,
         n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808,
         n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816,
         n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824,
         n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832,
         n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
         n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848,
         n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856,
         n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864,
         n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872,
         n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880,
         n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888,
         n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896,
         n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904,
         n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
         n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920,
         n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928,
         n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936,
         n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944,
         n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952,
         n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960,
         n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968,
         n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976,
         n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984,
         n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992,
         n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000,
         n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008,
         n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016,
         n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024,
         n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032,
         n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040,
         n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048,
         n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056,
         n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064,
         n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072,
         n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080,
         n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088,
         n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096,
         n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104,
         n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112,
         n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120,
         n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
         n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136,
         n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144,
         n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152,
         n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160,
         n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168,
         n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176,
         n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184,
         n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192,
         n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
         n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208,
         n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216,
         n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224,
         n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232,
         n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
         n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248,
         n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256,
         n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264,
         n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
         n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280,
         n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288,
         n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296,
         n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304,
         n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
         n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320,
         n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328,
         n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336,
         n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344,
         n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352,
         n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
         n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368,
         n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376,
         n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
         n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392,
         n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400,
         n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408,
         n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
         n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424,
         n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
         n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440,
         n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448,
         n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
         n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464,
         n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472,
         n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480,
         n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
         n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496,
         n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504,
         n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512,
         n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520,
         n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528,
         n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536,
         n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544,
         n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552,
         n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560,
         n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568,
         n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
         n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584,
         n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592,
         n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
         n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608,
         n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616,
         n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624,
         n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632,
         n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640,
         n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648,
         n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656,
         n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664,
         n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672,
         n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680,
         n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688,
         n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696,
         n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704,
         n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712,
         n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720,
         n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728,
         n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736,
         n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
         n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752,
         n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760,
         n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768,
         n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776,
         n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784,
         n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792,
         n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800,
         n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808,
         n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816,
         n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824,
         n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832,
         n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840,
         n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848,
         n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856,
         n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
         n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872,
         n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880,
         n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
         n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896,
         n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904,
         n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912,
         n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920,
         n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928,
         n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936,
         n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944,
         n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952,
         n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960,
         n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968,
         n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976,
         n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984,
         n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
         n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000,
         n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008,
         n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016,
         n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024,
         n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032,
         n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040,
         n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048,
         n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056,
         n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064,
         n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072,
         n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080,
         n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088,
         n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096,
         n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104,
         n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112,
         n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120,
         n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128,
         n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
         n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144,
         n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
         n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160,
         n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168,
         n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176,
         n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184,
         n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192,
         n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200,
         n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208,
         n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216,
         n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224,
         n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232,
         n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240,
         n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
         n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256,
         n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264,
         n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272,
         n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280,
         n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288,
         n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296,
         n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304,
         n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312,
         n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
         n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328,
         n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336,
         n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344,
         n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
         n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
         n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
         n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376,
         n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384,
         n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392,
         n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400,
         n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408,
         n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416,
         n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
         n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432,
         n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440,
         n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448,
         n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456,
         n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464,
         n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472,
         n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480,
         n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488,
         n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496,
         n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504,
         n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512,
         n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520,
         n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528,
         n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536,
         n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544,
         n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552,
         n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560,
         n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568,
         n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576,
         n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584,
         n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592,
         n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600,
         n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
         n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616,
         n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624,
         n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632,
         n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
         n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648,
         n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656,
         n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664,
         n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672,
         n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680,
         n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688,
         n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696,
         n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704,
         n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
         n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720,
         n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
         n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736,
         n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744,
         n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752,
         n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760,
         n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768,
         n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776,
         n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784,
         n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792,
         n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
         n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808,
         n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816,
         n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
         n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832,
         n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840,
         n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848,
         n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
         n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864,
         n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
         n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880,
         n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888,
         n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896,
         n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904,
         n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912,
         n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920,
         n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928,
         n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936,
         n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
         n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952,
         n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960,
         n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968,
         n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976,
         n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984,
         n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992,
         n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000,
         n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008,
         n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
         n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024,
         n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032,
         n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
         n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048,
         n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056,
         n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064,
         n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072,
         n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080,
         n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
         n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096,
         n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104,
         n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112,
         n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120,
         n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128,
         n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136,
         n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144,
         n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152,
         n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
         n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168,
         n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176,
         n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
         n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192,
         n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200,
         n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208,
         n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216,
         n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224,
         n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
         n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240,
         n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248,
         n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
         n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264,
         n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272,
         n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280,
         n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
         n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296,
         n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
         n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312,
         n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320,
         n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328,
         n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336,
         n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344,
         n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352,
         n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360,
         n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368,
         n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
         n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384,
         n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392,
         n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400,
         n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408,
         n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416,
         n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424,
         n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
         n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440,
         n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
         n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456,
         n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464,
         n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
         n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480,
         n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488,
         n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496,
         n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504,
         n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512,
         n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
         n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528,
         n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536,
         n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
         n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552,
         n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560,
         n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568,
         n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576,
         n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584,
         n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
         n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600,
         n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608,
         n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616,
         n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624,
         n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632,
         n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640,
         n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648,
         n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656,
         n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
         n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672,
         n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680,
         n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688,
         n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696,
         n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704,
         n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712,
         n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720,
         n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728,
         n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736,
         n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744,
         n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752,
         n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760,
         n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768,
         n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776,
         n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784,
         n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792,
         n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800,
         n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808,
         n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816,
         n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824,
         n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832,
         n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840,
         n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848,
         n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856,
         n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
         n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872,
         n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
         n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888,
         n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896,
         n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904,
         n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912,
         n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920,
         n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928,
         n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936,
         n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944,
         n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952,
         n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960,
         n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968,
         n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976,
         n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984,
         n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992,
         n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000,
         n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008,
         n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016,
         n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
         n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032,
         n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040,
         n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
         n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056,
         n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064,
         n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072,
         n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080,
         n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088,
         n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096,
         n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104,
         n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112,
         n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120,
         n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128,
         n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136,
         n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144,
         n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152,
         n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160,
         n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168,
         n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176,
         n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184,
         n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192,
         n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200,
         n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208,
         n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216,
         n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224,
         n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232,
         n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240,
         n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248,
         n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256,
         n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264,
         n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272,
         n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280,
         n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288,
         n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296,
         n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304,
         n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
         n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320,
         n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328,
         n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336,
         n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344,
         n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352,
         n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360,
         n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
         n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376,
         n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384,
         n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392,
         n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400,
         n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408,
         n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416,
         n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424,
         n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432,
         n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
         n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448,
         n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456,
         n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464,
         n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472,
         n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480,
         n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488,
         n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496,
         n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504,
         n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512,
         n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520,
         n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528,
         n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536,
         n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544,
         n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552,
         n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560,
         n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568,
         n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576,
         n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584,
         n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592,
         n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600,
         n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608,
         n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616,
         n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624,
         n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632,
         n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640,
         n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648,
         n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656,
         n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664,
         n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
         n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680,
         n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688,
         n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696,
         n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704,
         n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712,
         n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720,
         n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728,
         n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736,
         n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744,
         n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752,
         n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760,
         n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768,
         n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776,
         n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784,
         n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792,
         n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800,
         n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808,
         n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816,
         n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824,
         n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832,
         n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840,
         n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848,
         n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856,
         n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864,
         n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
         n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880,
         n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888,
         n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896,
         n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904,
         n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912,
         n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920,
         n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928,
         n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936,
         n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944,
         n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952,
         n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960,
         n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968,
         n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976,
         n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984,
         n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992,
         n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000,
         n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008,
         n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016,
         n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024,
         n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032,
         n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040,
         n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048,
         n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
         n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064,
         n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072,
         n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080,
         n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088,
         n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096,
         n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104,
         n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112,
         n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120,
         n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128,
         n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136,
         n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144,
         n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152,
         n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
         n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168,
         n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176,
         n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184,
         n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192,
         n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200,
         n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208,
         n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216,
         n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224,
         n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232,
         n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240,
         n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
         n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256,
         n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264,
         n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272,
         n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280,
         n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288,
         n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296,
         n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304,
         n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312,
         n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
         n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328,
         n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336,
         n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344,
         n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352,
         n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360,
         n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368,
         n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
         n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384,
         n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392,
         n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400,
         n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408,
         n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
         n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424,
         n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432,
         n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440,
         n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
         n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456,
         n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
         n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472,
         n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480,
         n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488,
         n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496,
         n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504,
         n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512,
         n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520,
         n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528,
         n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536,
         n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544,
         n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552,
         n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
         n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568,
         n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576,
         n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584,
         n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
         n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600,
         n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608,
         n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616,
         n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624,
         n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
         n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640,
         n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648,
         n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656,
         n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664,
         n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672,
         n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680,
         n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688,
         n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696,
         n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
         n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712,
         n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720,
         n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728,
         n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
         n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744,
         n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752,
         n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760,
         n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768,
         n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776,
         n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784,
         n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792,
         n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800,
         n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808,
         n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816,
         n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824,
         n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832,
         n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840,
         n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
         n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856,
         n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864,
         n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872,
         n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880,
         n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888,
         n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896,
         n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904,
         n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912,
         n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920,
         n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928,
         n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936,
         n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944,
         n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952,
         n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960,
         n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
         n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976,
         n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984,
         n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992,
         n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000,
         n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008,
         n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016,
         n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024,
         n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032,
         n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
         n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048,
         n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056,
         n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064,
         n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072,
         n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080,
         n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088,
         n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096,
         n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104,
         n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112,
         n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120,
         n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128,
         n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
         n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144,
         n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152,
         n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160,
         n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
         n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176,
         n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
         n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192,
         n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200,
         n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208,
         n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216,
         n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224,
         n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232,
         n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240,
         n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248,
         n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256,
         n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264,
         n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272,
         n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280,
         n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288,
         n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296,
         n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304,
         n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
         n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320,
         n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
         n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336,
         n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344,
         n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
         n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360,
         n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368,
         n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376,
         n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384,
         n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392,
         n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400,
         n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408,
         n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416,
         n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424,
         n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432,
         n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440,
         n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448,
         n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456,
         n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464,
         n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472,
         n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480,
         n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488,
         n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
         n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504,
         n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512,
         n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520,
         n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528,
         n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536,
         n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544,
         n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552,
         n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560,
         n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568,
         n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576,
         n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584,
         n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592,
         n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600,
         n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608,
         n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616,
         n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624,
         n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632,
         n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640,
         n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648,
         n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656,
         n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664,
         n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672,
         n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680,
         n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688,
         n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696,
         n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704,
         n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712,
         n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720,
         n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728,
         n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736,
         n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744,
         n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752,
         n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
         n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768,
         n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776,
         n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
         n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792,
         n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800,
         n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808,
         n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
         n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824,
         n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
         n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840,
         n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848,
         n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
         n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864,
         n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872,
         n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880,
         n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888,
         n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896,
         n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904,
         n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912,
         n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920,
         n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
         n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936,
         n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944,
         n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952,
         n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960,
         n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968,
         n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976,
         n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984,
         n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992,
         n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000,
         n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008,
         n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016,
         n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024,
         n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032,
         n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040,
         n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
         n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056,
         n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064,
         n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
         n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080,
         n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088,
         n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096,
         n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
         n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112,
         n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
         n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128,
         n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136,
         n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
         n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152,
         n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160,
         n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168,
         n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
         n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184,
         n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
         n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200,
         n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208,
         n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216,
         n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224,
         n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232,
         n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240,
         n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
         n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256,
         n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
         n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272,
         n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280,
         n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288,
         n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296,
         n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304,
         n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312,
         n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
         n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328,
         n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
         n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344,
         n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352,
         n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360,
         n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368,
         n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376,
         n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384,
         n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
         n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400,
         n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
         n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416,
         n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424,
         n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432,
         n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
         n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448,
         n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456,
         n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
         n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472,
         n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
         n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488,
         n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496,
         n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504,
         n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512,
         n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520,
         n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528,
         n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
         n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544,
         n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
         n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560,
         n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568,
         n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576,
         n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584,
         n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592,
         n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600,
         n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
         n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616,
         n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
         n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632,
         n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640,
         n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648,
         n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656,
         n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664,
         n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672,
         n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680,
         n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688,
         n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696,
         n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704,
         n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712,
         n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720,
         n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728,
         n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736,
         n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744,
         n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752,
         n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760,
         n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768,
         n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776,
         n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784,
         n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792,
         n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800,
         n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808,
         n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816,
         n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824,
         n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832,
         n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840,
         n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848,
         n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856,
         n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864,
         n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872,
         n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880,
         n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888,
         n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896,
         n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904,
         n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
         n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920,
         n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928,
         n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936,
         n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944,
         n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952,
         n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960,
         n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968,
         n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976,
         n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984,
         n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992,
         n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000,
         n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008,
         n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016,
         n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024,
         n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032,
         n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040,
         n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048,
         n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
         n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064,
         n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072,
         n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080,
         n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088,
         n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096,
         n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104,
         n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112,
         n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120,
         n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
         n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136,
         n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144,
         n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152,
         n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160,
         n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168,
         n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176,
         n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184,
         n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192,
         n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200,
         n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208,
         n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216,
         n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224,
         n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232,
         n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240,
         n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248,
         n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
         n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264,
         n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272,
         n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280,
         n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288,
         n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296,
         n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304,
         n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312,
         n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320,
         n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
         n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336,
         n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
         n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352,
         n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360,
         n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368,
         n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376,
         n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384,
         n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392,
         n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400,
         n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408,
         n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
         n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424,
         n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432,
         n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440,
         n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448,
         n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456,
         n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464,
         n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472,
         n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480,
         n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488,
         n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496,
         n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504,
         n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512,
         n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520,
         n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528,
         n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536,
         n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544,
         n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552,
         n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560,
         n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568,
         n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576,
         n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584,
         n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592,
         n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600,
         n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608,
         n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
         n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624,
         n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
         n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640,
         n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648,
         n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656,
         n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664,
         n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672,
         n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680,
         n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
         n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696,
         n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704,
         n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712,
         n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720,
         n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728,
         n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736,
         n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744,
         n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752,
         n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
         n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768,
         n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776,
         n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784,
         n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792,
         n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800,
         n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808,
         n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816,
         n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824,
         n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832,
         n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840,
         n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848,
         n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856,
         n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864,
         n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872,
         n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880,
         n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888,
         n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896,
         n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904,
         n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912,
         n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920,
         n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928,
         n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936,
         n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944,
         n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952,
         n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960,
         n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968,
         n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
         n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984,
         n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
         n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000,
         n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008,
         n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016,
         n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024,
         n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032,
         n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040,
         n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048,
         n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056,
         n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
         n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072,
         n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080,
         n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088,
         n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096,
         n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104,
         n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112,
         n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120,
         n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128,
         n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136,
         n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144,
         n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152,
         n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160,
         n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168,
         n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176,
         n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184,
         n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
         n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200,
         n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208,
         n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216,
         n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224,
         n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232,
         n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240,
         n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248,
         n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256,
         n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
         n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272,
         n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280,
         n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288,
         n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296,
         n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304,
         n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312,
         n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320,
         n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328,
         n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336,
         n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344,
         n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352,
         n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360,
         n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368,
         n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376,
         n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384,
         n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392,
         n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400,
         n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408,
         n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416,
         n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424,
         n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432,
         n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440,
         n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448,
         n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456,
         n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464,
         n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472,
         n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480,
         n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488,
         n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496,
         n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504,
         n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512,
         n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520,
         n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528,
         n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536,
         n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544,
         n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
         n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560,
         n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568,
         n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576,
         n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584,
         n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592,
         n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600,
         n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608,
         n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616,
         n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624,
         n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632,
         n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640,
         n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648,
         n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656,
         n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664,
         n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672,
         n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680,
         n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688,
         n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696,
         n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704,
         n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712,
         n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720,
         n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728,
         n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736,
         n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744,
         n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752,
         n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760,
         n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768,
         n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776,
         n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784,
         n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792,
         n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800,
         n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
         n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816,
         n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824,
         n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832,
         n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
         n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848,
         n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856,
         n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864,
         n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872,
         n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880,
         n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888,
         n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896,
         n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904,
         n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912,
         n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920,
         n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928,
         n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936,
         n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944,
         n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952,
         n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960,
         n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968,
         n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976,
         n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984,
         n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992,
         n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000,
         n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008,
         n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016,
         n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024,
         n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032,
         n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040,
         n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048,
         n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056,
         n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064,
         n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072,
         n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080,
         n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088,
         n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096,
         n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104,
         n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112,
         n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120,
         n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128,
         n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136,
         n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144,
         n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152,
         n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160,
         n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168,
         n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176,
         n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184,
         n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192,
         n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
         n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208,
         n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216,
         n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224,
         n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232,
         n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240,
         n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248,
         n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256,
         n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264,
         n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272,
         n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280,
         n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288,
         n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296,
         n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304,
         n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312,
         n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320,
         n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328,
         n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336,
         n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344,
         n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352,
         n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360,
         n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368,
         n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376,
         n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384,
         n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392,
         n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400,
         n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408,
         n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416,
         n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424,
         n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432,
         n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440,
         n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448,
         n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456,
         n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464,
         n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472,
         n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480,
         n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488,
         n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496,
         n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504,
         n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512,
         n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520,
         n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528,
         n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536,
         n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544,
         n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552,
         n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560,
         n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568,
         n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576,
         n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584,
         n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592,
         n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600,
         n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608,
         n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616,
         n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624,
         n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632,
         n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640,
         n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648,
         n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656,
         n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664,
         n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672,
         n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680,
         n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688,
         n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696,
         n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704,
         n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712,
         n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720,
         n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728,
         n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736,
         n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744,
         n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752,
         n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760,
         n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768,
         n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776,
         n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784,
         n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792,
         n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800,
         n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808,
         n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816,
         n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824,
         n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832,
         n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840,
         n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848,
         n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856,
         n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864,
         n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872,
         n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880,
         n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888,
         n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896,
         n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904,
         n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912,
         n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920,
         n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928,
         n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936,
         n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944,
         n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952,
         n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960,
         n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968,
         n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976,
         n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984,
         n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992,
         n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000,
         n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008,
         n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016,
         n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024,
         n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032,
         n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040,
         n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048,
         n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056,
         n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064,
         n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072,
         n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080,
         n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088,
         n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096,
         n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104,
         n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112,
         n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120,
         n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128,
         n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136,
         n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144,
         n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152,
         n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160,
         n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168,
         n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176,
         n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184,
         n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192,
         n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200,
         n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208,
         n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216,
         n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224,
         n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232,
         n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240,
         n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248,
         n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256,
         n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264,
         n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272,
         n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280,
         n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288,
         n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296,
         n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304,
         n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312,
         n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320,
         n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328,
         n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336,
         n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344,
         n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352,
         n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360,
         n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368,
         n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376,
         n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384,
         n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392,
         n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400,
         n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408,
         n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416,
         n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424,
         n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432,
         n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440,
         n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448,
         n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456,
         n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464,
         n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472,
         n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480,
         n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488,
         n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496,
         n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504,
         n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512,
         n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520,
         n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528,
         n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536,
         n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544,
         n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552,
         n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560,
         n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
         n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576,
         n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584,
         n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592,
         n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600,
         n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608,
         n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616,
         n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624,
         n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632,
         n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640,
         n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648,
         n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656,
         n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664,
         n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672,
         n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680,
         n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688,
         n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696,
         n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704,
         n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712,
         n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720,
         n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728,
         n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736,
         n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744,
         n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752,
         n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760,
         n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768,
         n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776,
         n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784,
         n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792,
         n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800,
         n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808,
         n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816,
         n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824,
         n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832,
         n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840,
         n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848,
         n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856,
         n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864,
         n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872,
         n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880,
         n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888,
         n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896,
         n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904,
         n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912,
         n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920,
         n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928,
         n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936,
         n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944,
         n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952,
         n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960,
         n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968,
         n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976,
         n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984,
         n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992,
         n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000,
         n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008,
         n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016,
         n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024,
         n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032,
         n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040,
         n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048,
         n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056,
         n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064,
         n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072,
         n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080,
         n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088,
         n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096,
         n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104,
         n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112,
         n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120,
         n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128,
         n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136,
         n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
         n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152,
         n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160,
         n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168,
         n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176,
         n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184,
         n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192,
         n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200,
         n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208,
         n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216,
         n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224,
         n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232,
         n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240,
         n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248,
         n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256,
         n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264,
         n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272,
         n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280,
         n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288,
         n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296,
         n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304,
         n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312,
         n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320,
         n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328,
         n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336,
         n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344,
         n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352,
         n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360,
         n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368,
         n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376,
         n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384,
         n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392,
         n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400,
         n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408,
         n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416,
         n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424,
         n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432,
         n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440,
         n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448,
         n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456,
         n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464,
         n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472,
         n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480,
         n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488,
         n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496,
         n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504,
         n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512,
         n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520,
         n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528,
         n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536,
         n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544,
         n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552,
         n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560,
         n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568,
         n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576,
         n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584,
         n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592,
         n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600,
         n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608,
         n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616,
         n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624,
         n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632,
         n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640,
         n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648,
         n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656,
         n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664,
         n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672,
         n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680,
         n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688,
         n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696,
         n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704,
         n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712,
         n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720,
         n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728,
         n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736,
         n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744,
         n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752,
         n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760,
         n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768,
         n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776,
         n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784,
         n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792,
         n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800,
         n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808,
         n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816,
         n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824,
         n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832,
         n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840,
         n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848,
         n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856,
         n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
         n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872,
         n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880,
         n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888,
         n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896,
         n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904,
         n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912,
         n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920,
         n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928,
         n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936,
         n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944,
         n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952,
         n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960,
         n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968,
         n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976,
         n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984,
         n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992,
         n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000,
         n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008,
         n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016,
         n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024,
         n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032,
         n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040,
         n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048,
         n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056,
         n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064,
         n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072,
         n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080,
         n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088,
         n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096,
         n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104,
         n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112,
         n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120,
         n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128,
         n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136,
         n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144,
         n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152,
         n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160,
         n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168,
         n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176,
         n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184,
         n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192,
         n56193, n56194, n56195;

  INV_X1 U23512 ( .A(1'b0), .ZN(n34468) );
  INV_X1 U23514 ( .A(1'b0), .ZN(n34467) );
  INV_X1 U23516 ( .A(1'b0), .ZN(n34466) );
  INV_X1 U23518 ( .A(1'b0), .ZN(n34465) );
  INV_X1 U23520 ( .A(1'b0), .ZN(n34464) );
  INV_X1 U23522 ( .A(1'b0), .ZN(n34461) );
  INV_X1 U23524 ( .A(1'b0), .ZN(n34460) );
  INV_X1 U23526 ( .A(1'b0), .ZN(n34459) );
  INV_X1 U23528 ( .A(1'b1), .ZN(n34458) );
  INV_X1 U23530 ( .A(1'b0), .ZN(n34457) );
  INV_X1 U23532 ( .A(1'b1), .ZN(n34423) );
  INV_X1 U23534 ( .A(1'b1), .ZN(n34422) );
  INV_X1 U23536 ( .A(1'b1), .ZN(n34421) );
  INV_X1 U23538 ( .A(1'b1), .ZN(n34420) );
  INV_X1 U23540 ( .A(1'b1), .ZN(n34419) );
  INV_X1 U23542 ( .A(1'b1), .ZN(n34418) );
  INV_X1 U23544 ( .A(1'b1), .ZN(n34417) );
  INV_X1 U23546 ( .A(1'b1), .ZN(n34416) );
  INV_X1 U23548 ( .A(1'b1), .ZN(n34415) );
  INV_X1 U23550 ( .A(1'b1), .ZN(n34414) );
  INV_X1 U23552 ( .A(1'b1), .ZN(n34413) );
  INV_X1 U23554 ( .A(1'b1), .ZN(n34412) );
  INV_X1 U23556 ( .A(1'b1), .ZN(n34411) );
  INV_X1 U23558 ( .A(1'b1), .ZN(n34410) );
  INV_X1 U23560 ( .A(1'b1), .ZN(n34409) );
  INV_X1 U23562 ( .A(1'b1), .ZN(n34408) );
  INV_X1 U23564 ( .A(1'b1), .ZN(n34407) );
  INV_X1 U23566 ( .A(1'b1), .ZN(n34406) );
  INV_X1 U23568 ( .A(1'b1), .ZN(n34405) );
  INV_X1 U23570 ( .A(1'b1), .ZN(n34404) );
  INV_X1 U23572 ( .A(1'b1), .ZN(n34403) );
  INV_X1 U23574 ( .A(1'b1), .ZN(n34402) );
  INV_X1 U23576 ( .A(1'b1), .ZN(n34401) );
  INV_X1 U23578 ( .A(1'b1), .ZN(n34400) );
  INV_X1 U23580 ( .A(1'b1), .ZN(n34399) );
  INV_X1 U23582 ( .A(1'b1), .ZN(n34398) );
  INV_X1 U23584 ( .A(1'b1), .ZN(n34397) );
  INV_X1 U23586 ( .A(1'b1), .ZN(n34396) );
  INV_X1 U23588 ( .A(1'b1), .ZN(n34395) );
  INV_X1 U23590 ( .A(1'b1), .ZN(n34394) );
  INV_X1 U23592 ( .A(1'b1), .ZN(n34393) );
  INV_X1 U23594 ( .A(1'b1), .ZN(n34392) );
  INV_X1 U23596 ( .A(1'b1), .ZN(n34391) );
  INV_X1 U23598 ( .A(1'b1), .ZN(n34390) );
  INV_X1 U23600 ( .A(1'b1), .ZN(n34389) );
  INV_X1 U23602 ( .A(1'b1), .ZN(n34388) );
  INV_X1 U23604 ( .A(1'b1), .ZN(n34387) );
  INV_X1 U23606 ( .A(1'b1), .ZN(n34386) );
  INV_X1 U23608 ( .A(1'b1), .ZN(n34385) );
  INV_X1 U23610 ( .A(1'b1), .ZN(n34384) );
  INV_X1 U23612 ( .A(1'b1), .ZN(n34383) );
  INV_X1 U23614 ( .A(1'b1), .ZN(n34382) );
  INV_X1 U23616 ( .A(1'b1), .ZN(n34381) );
  INV_X1 U23618 ( .A(1'b1), .ZN(n34380) );
  INV_X1 U23620 ( .A(1'b1), .ZN(n34379) );
  INV_X1 U23622 ( .A(1'b1), .ZN(n34378) );
  INV_X1 U23624 ( .A(1'b1), .ZN(n34377) );
  INV_X1 U23626 ( .A(1'b1), .ZN(n34376) );
  INV_X1 U23628 ( .A(1'b1), .ZN(n34375) );
  INV_X1 U23630 ( .A(1'b1), .ZN(n34374) );
  INV_X1 U23632 ( .A(1'b1), .ZN(n34373) );
  INV_X1 U23634 ( .A(1'b1), .ZN(n34372) );
  INV_X1 U23636 ( .A(1'b1), .ZN(n34371) );
  INV_X1 U23638 ( .A(1'b1), .ZN(n34370) );
  INV_X1 U23640 ( .A(1'b1), .ZN(n34369) );
  INV_X1 U23642 ( .A(1'b1), .ZN(n34368) );
  INV_X1 U23644 ( .A(1'b1), .ZN(n34367) );
  INV_X1 U23646 ( .A(1'b1), .ZN(n34366) );
  INV_X1 U23648 ( .A(1'b1), .ZN(n34365) );
  INV_X1 U23650 ( .A(1'b1), .ZN(n34364) );
  INV_X1 U23652 ( .A(1'b1), .ZN(n34363) );
  INV_X1 U23654 ( .A(1'b1), .ZN(n34362) );
  INV_X1 U23656 ( .A(1'b1), .ZN(n34361) );
  INV_X1 U23658 ( .A(1'b1), .ZN(n34360) );
  INV_X1 U23660 ( .A(1'b1), .ZN(n34359) );
  INV_X1 U23662 ( .A(1'b1), .ZN(n34358) );
  INV_X1 U23664 ( .A(1'b1), .ZN(n34357) );
  INV_X1 U23666 ( .A(1'b1), .ZN(n34356) );
  INV_X1 U23668 ( .A(1'b1), .ZN(n34355) );
  INV_X1 U23670 ( .A(1'b1), .ZN(n34354) );
  INV_X1 U23672 ( .A(1'b1), .ZN(n34353) );
  INV_X1 U23674 ( .A(1'b1), .ZN(n34352) );
  INV_X1 U23676 ( .A(1'b1), .ZN(n34351) );
  INV_X1 U23678 ( .A(1'b1), .ZN(n34350) );
  INV_X1 U23680 ( .A(1'b1), .ZN(n34349) );
  INV_X1 U23682 ( .A(1'b1), .ZN(n34348) );
  INV_X1 U23684 ( .A(1'b1), .ZN(n34347) );
  INV_X1 U23686 ( .A(1'b1), .ZN(n34346) );
  INV_X1 U23688 ( .A(1'b1), .ZN(n34345) );
  INV_X1 U23690 ( .A(1'b1), .ZN(n34344) );
  INV_X1 U23692 ( .A(1'b1), .ZN(n34343) );
  INV_X1 U23694 ( .A(1'b1), .ZN(n34342) );
  INV_X1 U23696 ( .A(1'b1), .ZN(n34341) );
  INV_X1 U23698 ( .A(1'b1), .ZN(n34340) );
  INV_X1 U23700 ( .A(1'b1), .ZN(n34339) );
  INV_X1 U23702 ( .A(1'b1), .ZN(n34338) );
  INV_X1 U23704 ( .A(1'b1), .ZN(n34337) );
  INV_X1 U23706 ( .A(1'b1), .ZN(n34336) );
  INV_X1 U23708 ( .A(1'b1), .ZN(n34335) );
  INV_X1 U23710 ( .A(1'b1), .ZN(n34334) );
  INV_X1 U23712 ( .A(1'b1), .ZN(n34333) );
  INV_X1 U23714 ( .A(1'b1), .ZN(n34332) );
  INV_X1 U23716 ( .A(1'b1), .ZN(n34331) );
  INV_X1 U23718 ( .A(1'b1), .ZN(n34330) );
  INV_X1 U23720 ( .A(1'b1), .ZN(n34329) );
  INV_X1 U23722 ( .A(1'b1), .ZN(n34328) );
  INV_X1 U23724 ( .A(1'b1), .ZN(n34327) );
  INV_X1 U23726 ( .A(1'b1), .ZN(n34326) );
  INV_X1 U23728 ( .A(1'b1), .ZN(n34325) );
  INV_X1 U23730 ( .A(1'b1), .ZN(n34324) );
  INV_X1 U23732 ( .A(1'b1), .ZN(n34323) );
  INV_X1 U23734 ( .A(1'b1), .ZN(n34322) );
  INV_X1 U23736 ( .A(1'b1), .ZN(n34321) );
  INV_X1 U23738 ( .A(1'b1), .ZN(n34320) );
  INV_X1 U23740 ( .A(1'b1), .ZN(n34319) );
  INV_X1 U23742 ( .A(1'b1), .ZN(n34318) );
  INV_X1 U23744 ( .A(1'b1), .ZN(n34317) );
  INV_X1 U23746 ( .A(1'b1), .ZN(n34316) );
  INV_X1 U23748 ( .A(1'b1), .ZN(n34315) );
  INV_X1 U23750 ( .A(1'b1), .ZN(n34314) );
  INV_X1 U23752 ( .A(1'b1), .ZN(n34313) );
  INV_X1 U23754 ( .A(1'b1), .ZN(n34312) );
  INV_X1 U23756 ( .A(1'b1), .ZN(n34311) );
  INV_X1 U23758 ( .A(1'b1), .ZN(n34310) );
  INV_X1 U23760 ( .A(1'b1), .ZN(n34309) );
  INV_X1 U23762 ( .A(1'b1), .ZN(n34308) );
  INV_X1 U23764 ( .A(1'b1), .ZN(n34307) );
  INV_X1 U23766 ( .A(1'b1), .ZN(n34306) );
  INV_X1 U23768 ( .A(1'b1), .ZN(n34305) );
  INV_X1 U23770 ( .A(1'b1), .ZN(n34304) );
  INV_X1 U23772 ( .A(1'b1), .ZN(n34303) );
  INV_X1 U23774 ( .A(1'b1), .ZN(n34302) );
  INV_X1 U23776 ( .A(1'b1), .ZN(n34301) );
  INV_X1 U23778 ( .A(1'b1), .ZN(n34300) );
  INV_X1 U23780 ( .A(1'b1), .ZN(n34299) );
  INV_X1 U23782 ( .A(1'b1), .ZN(n34298) );
  INV_X1 U23784 ( .A(1'b1), .ZN(n34297) );
  INV_X1 U23786 ( .A(1'b1), .ZN(n34296) );
  INV_X1 U23788 ( .A(1'b1), .ZN(n34295) );
  INV_X1 U23790 ( .A(1'b1), .ZN(n34294) );
  INV_X1 U23792 ( .A(1'b1), .ZN(n34293) );
  INV_X1 U23794 ( .A(1'b1), .ZN(n34292) );
  INV_X1 U23796 ( .A(1'b1), .ZN(n34291) );
  INV_X1 U23798 ( .A(1'b1), .ZN(n34290) );
  INV_X1 U23800 ( .A(1'b1), .ZN(n34289) );
  INV_X1 U23802 ( .A(1'b1), .ZN(n34288) );
  INV_X1 U23804 ( .A(1'b1), .ZN(n34287) );
  INV_X1 U23806 ( .A(1'b1), .ZN(n34286) );
  INV_X1 U23808 ( .A(1'b1), .ZN(n34285) );
  INV_X1 U23810 ( .A(1'b1), .ZN(n34284) );
  INV_X1 U23812 ( .A(1'b1), .ZN(n34283) );
  INV_X1 U23814 ( .A(1'b1), .ZN(n34282) );
  INV_X1 U23816 ( .A(1'b1), .ZN(n34281) );
  INV_X1 U23818 ( .A(1'b1), .ZN(n34280) );
  INV_X1 U23820 ( .A(1'b1), .ZN(n34279) );
  INV_X1 U23822 ( .A(1'b1), .ZN(n34278) );
  INV_X1 U23824 ( .A(1'b1), .ZN(n34277) );
  INV_X1 U23826 ( .A(1'b1), .ZN(n34276) );
  INV_X1 U23828 ( .A(1'b1), .ZN(n34275) );
  INV_X1 U23830 ( .A(1'b1), .ZN(n34274) );
  INV_X1 U23832 ( .A(1'b1), .ZN(n34273) );
  INV_X1 U23834 ( .A(1'b1), .ZN(n34272) );
  INV_X1 U23836 ( .A(1'b1), .ZN(n34271) );
  INV_X1 U23838 ( .A(1'b1), .ZN(n34270) );
  INV_X1 U23840 ( .A(1'b1), .ZN(n34269) );
  INV_X1 U23842 ( .A(1'b1), .ZN(n34268) );
  INV_X1 U23844 ( .A(1'b1), .ZN(n34267) );
  INV_X1 U23846 ( .A(1'b1), .ZN(n34266) );
  INV_X1 U23848 ( .A(1'b1), .ZN(n34265) );
  INV_X1 U23850 ( .A(1'b1), .ZN(n34264) );
  INV_X1 U23852 ( .A(1'b1), .ZN(n34263) );
  INV_X1 U23854 ( .A(1'b1), .ZN(n34262) );
  INV_X1 U23856 ( .A(1'b1), .ZN(n34261) );
  INV_X1 U23858 ( .A(1'b1), .ZN(n34260) );
  INV_X1 U23860 ( .A(1'b1), .ZN(n34259) );
  INV_X1 U23862 ( .A(1'b1), .ZN(n34258) );
  INV_X1 U23864 ( .A(1'b1), .ZN(n34257) );
  INV_X1 U23866 ( .A(1'b1), .ZN(n34256) );
  INV_X1 U23868 ( .A(1'b1), .ZN(n34255) );
  INV_X1 U23870 ( .A(1'b1), .ZN(n34254) );
  INV_X1 U23872 ( .A(1'b1), .ZN(n34253) );
  INV_X1 U23874 ( .A(1'b1), .ZN(n34252) );
  INV_X1 U23876 ( .A(1'b1), .ZN(n34251) );
  INV_X1 U23878 ( .A(1'b1), .ZN(n34250) );
  INV_X1 U23880 ( .A(1'b1), .ZN(n34249) );
  INV_X1 U23882 ( .A(1'b1), .ZN(n34248) );
  INV_X1 U23884 ( .A(1'b1), .ZN(n34247) );
  INV_X1 U23886 ( .A(1'b1), .ZN(n34246) );
  INV_X1 U23888 ( .A(1'b1), .ZN(n34245) );
  INV_X1 U23890 ( .A(1'b1), .ZN(n34244) );
  INV_X1 U23892 ( .A(1'b1), .ZN(n34243) );
  INV_X1 U23894 ( .A(1'b1), .ZN(n34242) );
  INV_X1 U23896 ( .A(1'b1), .ZN(n34241) );
  INV_X1 U23898 ( .A(1'b1), .ZN(n34240) );
  INV_X1 U23900 ( .A(1'b1), .ZN(n34239) );
  INV_X1 U23902 ( .A(1'b1), .ZN(n34238) );
  INV_X1 U23904 ( .A(1'b1), .ZN(n34237) );
  INV_X1 U23906 ( .A(1'b1), .ZN(n34236) );
  INV_X1 U23908 ( .A(1'b1), .ZN(n34235) );
  INV_X1 U23910 ( .A(1'b1), .ZN(n34234) );
  INV_X1 U23912 ( .A(1'b1), .ZN(n34233) );
  INV_X1 U23914 ( .A(1'b1), .ZN(n34232) );
  INV_X1 U23916 ( .A(1'b1), .ZN(n34231) );
  INV_X1 U23918 ( .A(1'b1), .ZN(n34230) );
  INV_X1 U23920 ( .A(1'b1), .ZN(n34229) );
  INV_X1 U23922 ( .A(1'b1), .ZN(n34228) );
  INV_X1 U23924 ( .A(1'b1), .ZN(n34227) );
  INV_X1 U23926 ( .A(1'b1), .ZN(n34226) );
  INV_X1 U23928 ( .A(1'b1), .ZN(n34225) );
  INV_X1 U23930 ( .A(1'b1), .ZN(n34224) );
  INV_X1 U23932 ( .A(1'b1), .ZN(n34223) );
  INV_X1 U23934 ( .A(1'b1), .ZN(n34222) );
  INV_X1 U23936 ( .A(1'b1), .ZN(n34221) );
  INV_X1 U23938 ( .A(1'b1), .ZN(n34220) );
  INV_X1 U23940 ( .A(1'b1), .ZN(n34219) );
  INV_X1 U23942 ( .A(1'b1), .ZN(n34218) );
  INV_X1 U23944 ( .A(1'b1), .ZN(n34217) );
  INV_X1 U23946 ( .A(1'b1), .ZN(n34216) );
  INV_X1 U23948 ( .A(1'b1), .ZN(n34215) );
  INV_X1 U23950 ( .A(1'b1), .ZN(n34214) );
  INV_X1 U23952 ( .A(1'b1), .ZN(n34213) );
  INV_X1 U23954 ( .A(1'b1), .ZN(n34212) );
  INV_X1 U23956 ( .A(1'b1), .ZN(n34211) );
  INV_X1 U23958 ( .A(1'b1), .ZN(n34210) );
  INV_X1 U23960 ( .A(1'b1), .ZN(n34209) );
  INV_X1 U23962 ( .A(1'b1), .ZN(n34208) );
  INV_X1 U23964 ( .A(1'b1), .ZN(n34207) );
  INV_X1 U23966 ( .A(1'b1), .ZN(n34206) );
  INV_X1 U23968 ( .A(1'b1), .ZN(n34205) );
  INV_X1 U23970 ( .A(1'b1), .ZN(n34204) );
  INV_X1 U23972 ( .A(1'b1), .ZN(n34203) );
  INV_X1 U23974 ( .A(1'b1), .ZN(n34202) );
  INV_X1 U23976 ( .A(1'b1), .ZN(n34201) );
  INV_X1 U23978 ( .A(1'b1), .ZN(n34200) );
  INV_X1 U23980 ( .A(1'b1), .ZN(n34199) );
  INV_X1 U23982 ( .A(1'b1), .ZN(n34198) );
  INV_X1 U23984 ( .A(1'b1), .ZN(n34197) );
  INV_X1 U23986 ( .A(1'b1), .ZN(n34196) );
  INV_X1 U23988 ( .A(1'b1), .ZN(n34195) );
  INV_X1 U23990 ( .A(1'b1), .ZN(n34194) );
  INV_X1 U23992 ( .A(1'b1), .ZN(n34193) );
  INV_X1 U23994 ( .A(1'b1), .ZN(n34192) );
  INV_X1 U23996 ( .A(1'b1), .ZN(n34191) );
  INV_X1 U23998 ( .A(1'b1), .ZN(n34190) );
  INV_X1 U24000 ( .A(1'b1), .ZN(n34189) );
  INV_X1 U24002 ( .A(1'b1), .ZN(n34188) );
  INV_X1 U24004 ( .A(1'b1), .ZN(n34187) );
  INV_X1 U24006 ( .A(1'b1), .ZN(n34186) );
  INV_X1 U24008 ( .A(1'b1), .ZN(n34185) );
  INV_X1 U24010 ( .A(1'b1), .ZN(n34184) );
  INV_X1 U24012 ( .A(1'b1), .ZN(n34183) );
  INV_X1 U24014 ( .A(1'b1), .ZN(n34182) );
  INV_X1 U24016 ( .A(1'b1), .ZN(n34181) );
  INV_X1 U24018 ( .A(1'b1), .ZN(n34180) );
  INV_X1 U24020 ( .A(1'b1), .ZN(n34179) );
  INV_X1 U24022 ( .A(1'b1), .ZN(n34178) );
  INV_X1 U24024 ( .A(1'b1), .ZN(n34177) );
  INV_X1 U24026 ( .A(1'b1), .ZN(n34176) );
  INV_X1 U24028 ( .A(1'b1), .ZN(n34175) );
  INV_X1 U24030 ( .A(1'b1), .ZN(n34174) );
  INV_X1 U24032 ( .A(1'b1), .ZN(n34173) );
  INV_X1 U24034 ( .A(1'b1), .ZN(n34172) );
  INV_X1 U24036 ( .A(1'b1), .ZN(n34171) );
  INV_X1 U24038 ( .A(1'b1), .ZN(n34170) );
  INV_X1 U24040 ( .A(1'b1), .ZN(n34169) );
  INV_X1 U24042 ( .A(1'b1), .ZN(n34168) );
  INV_X1 U24044 ( .A(1'b1), .ZN(n34167) );
  INV_X1 U24046 ( .A(1'b1), .ZN(n34166) );
  INV_X1 U24048 ( .A(1'b1), .ZN(n34165) );
  INV_X1 U24050 ( .A(1'b1), .ZN(n34164) );
  INV_X1 U24052 ( .A(1'b1), .ZN(n34163) );
  INV_X1 U24054 ( .A(1'b1), .ZN(n34162) );
  INV_X1 U24056 ( .A(1'b1), .ZN(n34161) );
  INV_X1 U24058 ( .A(1'b1), .ZN(n34160) );
  INV_X1 U24060 ( .A(1'b1), .ZN(n34159) );
  INV_X1 U24062 ( .A(1'b1), .ZN(n34158) );
  INV_X1 U24064 ( .A(1'b1), .ZN(n34157) );
  INV_X1 U24066 ( .A(1'b1), .ZN(n34156) );
  INV_X1 U24068 ( .A(1'b1), .ZN(n34155) );
  INV_X1 U24070 ( .A(1'b1), .ZN(n34154) );
  INV_X1 U24072 ( .A(1'b1), .ZN(n34153) );
  INV_X1 U24074 ( .A(1'b1), .ZN(n34152) );
  INV_X1 U24076 ( .A(1'b1), .ZN(n34151) );
  INV_X1 U24078 ( .A(1'b1), .ZN(n34150) );
  INV_X1 U24080 ( .A(1'b1), .ZN(n34149) );
  INV_X1 U24082 ( .A(1'b1), .ZN(n34148) );
  INV_X1 U24084 ( .A(1'b1), .ZN(n34147) );
  INV_X1 U24086 ( .A(1'b1), .ZN(n34146) );
  INV_X1 U24088 ( .A(1'b1), .ZN(n34145) );
  INV_X1 U24090 ( .A(1'b1), .ZN(n34144) );
  INV_X1 U24092 ( .A(1'b1), .ZN(n34143) );
  INV_X1 U24094 ( .A(1'b1), .ZN(n34142) );
  INV_X1 U24096 ( .A(1'b1), .ZN(n34141) );
  INV_X1 U24098 ( .A(1'b1), .ZN(n34140) );
  INV_X1 U24100 ( .A(1'b1), .ZN(n34139) );
  INV_X1 U24102 ( .A(1'b1), .ZN(n34138) );
  INV_X1 U24104 ( .A(1'b1), .ZN(n34137) );
  INV_X1 U24106 ( .A(1'b1), .ZN(n34136) );
  INV_X1 U24108 ( .A(1'b1), .ZN(n34135) );
  INV_X1 U24110 ( .A(1'b1), .ZN(n34134) );
  INV_X1 U24112 ( .A(1'b1), .ZN(n34133) );
  INV_X1 U24114 ( .A(1'b1), .ZN(n34132) );
  INV_X1 U24116 ( .A(1'b1), .ZN(n34131) );
  INV_X1 U24118 ( .A(1'b1), .ZN(n34130) );
  INV_X1 U24120 ( .A(1'b1), .ZN(n34129) );
  INV_X1 U24122 ( .A(1'b1), .ZN(n34128) );
  INV_X1 U24124 ( .A(1'b1), .ZN(n34127) );
  INV_X1 U24126 ( .A(1'b1), .ZN(n34126) );
  INV_X1 U24128 ( .A(1'b1), .ZN(n34125) );
  INV_X1 U24130 ( .A(1'b1), .ZN(n34124) );
  INV_X1 U24132 ( .A(1'b1), .ZN(n34123) );
  INV_X1 U24134 ( .A(1'b1), .ZN(n34122) );
  INV_X1 U24136 ( .A(1'b1), .ZN(n34121) );
  INV_X1 U24138 ( .A(1'b1), .ZN(n34120) );
  INV_X1 U24140 ( .A(1'b1), .ZN(n34119) );
  INV_X1 U24142 ( .A(1'b1), .ZN(n34118) );
  INV_X1 U24144 ( .A(1'b1), .ZN(n34117) );
  INV_X1 U24146 ( .A(1'b1), .ZN(n34116) );
  INV_X1 U24148 ( .A(1'b1), .ZN(n34115) );
  INV_X1 U24150 ( .A(1'b1), .ZN(n34114) );
  INV_X1 U24152 ( .A(1'b1), .ZN(n34113) );
  INV_X1 U24154 ( .A(1'b1), .ZN(n34112) );
  INV_X1 U24156 ( .A(1'b1), .ZN(n34111) );
  INV_X1 U24158 ( .A(1'b1), .ZN(n34110) );
  INV_X1 U24160 ( .A(1'b1), .ZN(n34109) );
  INV_X1 U24162 ( .A(1'b1), .ZN(n34108) );
  INV_X1 U24164 ( .A(1'b1), .ZN(n34107) );
  INV_X1 U24166 ( .A(1'b1), .ZN(n34106) );
  INV_X1 U24168 ( .A(1'b1), .ZN(n34105) );
  INV_X1 U24170 ( .A(1'b1), .ZN(n34104) );
  INV_X1 U24172 ( .A(1'b1), .ZN(n34103) );
  INV_X1 U24174 ( .A(1'b1), .ZN(n34102) );
  INV_X1 U24176 ( .A(1'b1), .ZN(n34101) );
  INV_X1 U24178 ( .A(1'b1), .ZN(n34100) );
  INV_X1 U24180 ( .A(1'b1), .ZN(n34099) );
  INV_X1 U24182 ( .A(1'b1), .ZN(n34098) );
  INV_X1 U24184 ( .A(1'b1), .ZN(n34097) );
  INV_X1 U24186 ( .A(1'b1), .ZN(n34096) );
  INV_X1 U24188 ( .A(1'b1), .ZN(n34095) );
  INV_X1 U24190 ( .A(1'b1), .ZN(n34094) );
  INV_X1 U24192 ( .A(1'b1), .ZN(n34093) );
  INV_X1 U24194 ( .A(1'b1), .ZN(n34092) );
  INV_X1 U24196 ( .A(1'b1), .ZN(n34091) );
  INV_X1 U24198 ( .A(1'b1), .ZN(n34090) );
  INV_X1 U24200 ( .A(1'b1), .ZN(n34089) );
  INV_X1 U24202 ( .A(1'b1), .ZN(n34088) );
  INV_X1 U24204 ( .A(1'b1), .ZN(n34087) );
  INV_X1 U24206 ( .A(1'b1), .ZN(n34086) );
  INV_X1 U24208 ( .A(1'b1), .ZN(n34085) );
  INV_X1 U24210 ( .A(1'b1), .ZN(n34084) );
  INV_X1 U24212 ( .A(1'b1), .ZN(n34083) );
  INV_X1 U24214 ( .A(1'b1), .ZN(n34082) );
  INV_X1 U24216 ( .A(1'b1), .ZN(n34081) );
  INV_X1 U24218 ( .A(1'b1), .ZN(n34080) );
  INV_X1 U24220 ( .A(1'b1), .ZN(n34079) );
  INV_X1 U24222 ( .A(1'b1), .ZN(n34078) );
  INV_X1 U24224 ( .A(1'b1), .ZN(n34077) );
  INV_X1 U24226 ( .A(1'b1), .ZN(n34076) );
  INV_X1 U24228 ( .A(1'b1), .ZN(n34075) );
  INV_X1 U24230 ( .A(1'b1), .ZN(n34074) );
  INV_X1 U24232 ( .A(1'b1), .ZN(n34073) );
  INV_X1 U24234 ( .A(1'b1), .ZN(n34072) );
  INV_X1 U24236 ( .A(1'b1), .ZN(n34071) );
  INV_X1 U24238 ( .A(1'b1), .ZN(n34070) );
  INV_X1 U24240 ( .A(1'b1), .ZN(n34069) );
  INV_X1 U24242 ( .A(1'b1), .ZN(n34068) );
  INV_X1 U24244 ( .A(1'b1), .ZN(n34067) );
  INV_X1 U24246 ( .A(1'b1), .ZN(n34066) );
  INV_X1 U24248 ( .A(1'b1), .ZN(n34065) );
  INV_X1 U24250 ( .A(1'b1), .ZN(n34064) );
  INV_X1 U24252 ( .A(1'b1), .ZN(n34063) );
  INV_X1 U24254 ( .A(1'b1), .ZN(n34062) );
  INV_X1 U24256 ( .A(1'b1), .ZN(n34061) );
  INV_X1 U24258 ( .A(1'b1), .ZN(n34060) );
  INV_X1 U24260 ( .A(1'b1), .ZN(n34059) );
  INV_X1 U24262 ( .A(1'b1), .ZN(n34058) );
  INV_X1 U24264 ( .A(1'b1), .ZN(n34057) );
  INV_X1 U24266 ( .A(1'b1), .ZN(n34056) );
  INV_X1 U24268 ( .A(1'b1), .ZN(n34055) );
  INV_X1 U24270 ( .A(1'b1), .ZN(n34054) );
  INV_X1 U24272 ( .A(1'b1), .ZN(n34053) );
  INV_X1 U24274 ( .A(1'b1), .ZN(n34052) );
  INV_X1 U24276 ( .A(1'b1), .ZN(n34051) );
  INV_X1 U24278 ( .A(1'b1), .ZN(n34050) );
  INV_X1 U24280 ( .A(1'b1), .ZN(n34049) );
  INV_X1 U24282 ( .A(1'b1), .ZN(n34048) );
  INV_X1 U24284 ( .A(1'b1), .ZN(n34047) );
  INV_X1 U24286 ( .A(1'b1), .ZN(n34046) );
  INV_X1 U24288 ( .A(1'b1), .ZN(n34045) );
  INV_X1 U24290 ( .A(1'b1), .ZN(n34044) );
  INV_X1 U24292 ( .A(1'b1), .ZN(n34043) );
  INV_X1 U24294 ( .A(1'b1), .ZN(n34042) );
  INV_X1 U24296 ( .A(1'b1), .ZN(n34041) );
  INV_X1 U24298 ( .A(1'b1), .ZN(n34040) );
  INV_X1 U24300 ( .A(1'b1), .ZN(n34039) );
  INV_X1 U24302 ( .A(1'b1), .ZN(n34038) );
  INV_X1 U24304 ( .A(1'b1), .ZN(n34037) );
  INV_X1 U24306 ( .A(1'b1), .ZN(n34036) );
  INV_X1 U24308 ( .A(1'b1), .ZN(n34035) );
  INV_X1 U24310 ( .A(1'b1), .ZN(n34034) );
  INV_X1 U24312 ( .A(1'b1), .ZN(n34033) );
  INV_X1 U24314 ( .A(1'b1), .ZN(n34032) );
  INV_X1 U24316 ( .A(1'b1), .ZN(n34031) );
  INV_X1 U24318 ( .A(1'b1), .ZN(n34030) );
  INV_X1 U24320 ( .A(1'b1), .ZN(n34029) );
  INV_X1 U24322 ( .A(1'b1), .ZN(n34028) );
  INV_X1 U24324 ( .A(1'b1), .ZN(n34027) );
  INV_X1 U24326 ( .A(1'b1), .ZN(n34026) );
  INV_X1 U24328 ( .A(1'b1), .ZN(n34025) );
  INV_X1 U24330 ( .A(1'b1), .ZN(n34024) );
  INV_X1 U24332 ( .A(1'b1), .ZN(n34023) );
  INV_X1 U24334 ( .A(1'b1), .ZN(n34022) );
  INV_X1 U24336 ( .A(1'b1), .ZN(n34021) );
  INV_X1 U24338 ( .A(1'b1), .ZN(n34020) );
  INV_X1 U24340 ( .A(1'b1), .ZN(n34019) );
  INV_X1 U24342 ( .A(1'b1), .ZN(n34018) );
  INV_X1 U24344 ( .A(1'b1), .ZN(n34017) );
  INV_X1 U24346 ( .A(1'b1), .ZN(n34016) );
  INV_X1 U24348 ( .A(1'b1), .ZN(n34015) );
  INV_X1 U24350 ( .A(1'b1), .ZN(n34014) );
  INV_X1 U24352 ( .A(1'b1), .ZN(n34013) );
  INV_X1 U24354 ( .A(1'b1), .ZN(n34012) );
  INV_X1 U24356 ( .A(1'b1), .ZN(n34011) );
  INV_X1 U24358 ( .A(1'b1), .ZN(n34010) );
  INV_X1 U24360 ( .A(1'b1), .ZN(n34009) );
  INV_X1 U24362 ( .A(1'b1), .ZN(n34008) );
  INV_X1 U24364 ( .A(1'b1), .ZN(n34007) );
  INV_X1 U24366 ( .A(1'b1), .ZN(n34006) );
  INV_X1 U24368 ( .A(1'b1), .ZN(n34005) );
  INV_X1 U24370 ( .A(1'b1), .ZN(n34004) );
  INV_X1 U24372 ( .A(1'b1), .ZN(n34003) );
  INV_X1 U24374 ( .A(1'b1), .ZN(n34002) );
  INV_X1 U24376 ( .A(1'b1), .ZN(n34001) );
  INV_X1 U24378 ( .A(1'b1), .ZN(n34000) );
  INV_X1 U24380 ( .A(1'b1), .ZN(n33999) );
  INV_X1 U24382 ( .A(1'b1), .ZN(n33998) );
  INV_X1 U24384 ( .A(1'b1), .ZN(n33997) );
  INV_X1 U24386 ( .A(1'b1), .ZN(n33996) );
  INV_X1 U24388 ( .A(1'b1), .ZN(n33995) );
  INV_X1 U24390 ( .A(1'b1), .ZN(n33994) );
  INV_X1 U24392 ( .A(1'b1), .ZN(n33993) );
  INV_X1 U24394 ( .A(1'b1), .ZN(n33992) );
  INV_X1 U24396 ( .A(1'b1), .ZN(n33991) );
  INV_X1 U24398 ( .A(1'b1), .ZN(n33990) );
  INV_X1 U24400 ( .A(1'b1), .ZN(n33989) );
  INV_X1 U24402 ( .A(1'b1), .ZN(n33988) );
  INV_X1 U24404 ( .A(1'b1), .ZN(n33987) );
  INV_X1 U24406 ( .A(1'b1), .ZN(n33986) );
  INV_X1 U24408 ( .A(1'b1), .ZN(n33985) );
  INV_X1 U24410 ( .A(1'b1), .ZN(n33984) );
  INV_X1 U24412 ( .A(1'b1), .ZN(n33983) );
  INV_X1 U24414 ( .A(1'b1), .ZN(n33982) );
  INV_X1 U24416 ( .A(1'b1), .ZN(n33981) );
  INV_X1 U24418 ( .A(1'b1), .ZN(n33980) );
  INV_X1 U24420 ( .A(1'b1), .ZN(n33979) );
  INV_X1 U24422 ( .A(1'b1), .ZN(n33978) );
  INV_X1 U24424 ( .A(1'b1), .ZN(n33977) );
  INV_X1 U24426 ( .A(1'b1), .ZN(n33976) );
  INV_X1 U24428 ( .A(1'b1), .ZN(n33975) );
  INV_X1 U24430 ( .A(1'b1), .ZN(n33974) );
  INV_X1 U24432 ( .A(1'b1), .ZN(n33973) );
  INV_X1 U24434 ( .A(1'b1), .ZN(n33972) );
  INV_X1 U24436 ( .A(1'b1), .ZN(n33971) );
  INV_X1 U24438 ( .A(1'b1), .ZN(n33970) );
  INV_X1 U24440 ( .A(1'b1), .ZN(n33969) );
  INV_X1 U24442 ( .A(1'b1), .ZN(n33968) );
  INV_X1 U24444 ( .A(1'b1), .ZN(n33967) );
  INV_X1 U24446 ( .A(1'b1), .ZN(n33966) );
  INV_X1 U24448 ( .A(1'b1), .ZN(n33965) );
  INV_X1 U24450 ( .A(1'b1), .ZN(n33964) );
  INV_X1 U24452 ( .A(1'b1), .ZN(n33963) );
  INV_X1 U24454 ( .A(1'b1), .ZN(n33962) );
  INV_X1 U24456 ( .A(1'b1), .ZN(n33961) );
  INV_X1 U24458 ( .A(1'b1), .ZN(n33960) );
  INV_X1 U24460 ( .A(1'b1), .ZN(n33959) );
  INV_X1 U24462 ( .A(1'b1), .ZN(n33958) );
  INV_X1 U24464 ( .A(1'b1), .ZN(n33957) );
  INV_X1 U24466 ( .A(1'b1), .ZN(n33956) );
  INV_X1 U24468 ( .A(1'b1), .ZN(n33955) );
  INV_X1 U24470 ( .A(1'b1), .ZN(n33954) );
  INV_X1 U24472 ( .A(1'b1), .ZN(n33953) );
  INV_X1 U24474 ( .A(1'b1), .ZN(n33952) );
  INV_X1 U24476 ( .A(1'b1), .ZN(n33951) );
  INV_X1 U24478 ( .A(1'b1), .ZN(n33950) );
  INV_X1 U24480 ( .A(1'b1), .ZN(n33949) );
  INV_X1 U24482 ( .A(1'b1), .ZN(n33948) );
  INV_X1 U24484 ( .A(1'b1), .ZN(n33947) );
  INV_X1 U24486 ( .A(1'b1), .ZN(n33946) );
  INV_X1 U24488 ( .A(1'b1), .ZN(n33945) );
  INV_X1 U24490 ( .A(1'b1), .ZN(n33944) );
  INV_X1 U24492 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N654) );
  INV_X1 U24494 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N653) );
  INV_X1 U24496 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N652) );
  INV_X1 U24498 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N651) );
  INV_X1 U24500 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N650) );
  INV_X1 U24502 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N649) );
  INV_X1 U24504 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N648) );
  INV_X1 U24506 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N647) );
  INV_X1 U24508 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N646) );
  INV_X1 U24510 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N645) );
  INV_X1 U24512 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N644) );
  INV_X1 U24514 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N643) );
  INV_X1 U24516 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N642) );
  INV_X1 U24518 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N641) );
  INV_X1 U24520 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N640) );
  INV_X1 U24522 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N639) );
  INV_X1 U24524 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N638) );
  INV_X1 U24526 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N637) );
  INV_X1 U24528 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N636) );
  INV_X1 U24530 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N635) );
  INV_X1 U24532 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N634) );
  INV_X1 U24534 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N633) );
  INV_X1 U24536 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N632) );
  INV_X1 U24538 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N631) );
  INV_X1 U24540 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N630) );
  INV_X1 U24542 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N629) );
  INV_X1 U24544 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N628) );
  INV_X1 U24546 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N627) );
  INV_X1 U24548 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N626) );
  INV_X1 U24550 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N625) );
  INV_X1 U24552 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N624) );
  INV_X1 U24554 ( .A(1'b1), .ZN(p_wishbone_rx_fifo_N623) );
  INV_X1 U24556 ( .A(1'b1), .ZN(p_rxethmac1_crcrx_N3) );
  INV_X1 U24558 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N7) );
  INV_X1 U24560 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N11) );
  INV_X1 U24562 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N12) );
  INV_X1 U24564 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N10) );
  INV_X1 U24566 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N8) );
  INV_X1 U24568 ( .A(1'b1), .ZN(p_rxethmac1_crcrx_N5) );
  INV_X1 U24570 ( .A(1'b0), .ZN(p_rxethmac1_crcrx_N13) );
  INV_X1 U24572 ( .A(1'b0), .ZN(n35881) );
  INV_X1 U24574 ( .A(1'b0), .ZN(n35880) );
  INV_X1 U24576 ( .A(1'b0), .ZN(n35879) );
  INV_X1 U24578 ( .A(1'b0), .ZN(n35878) );
  INV_X1 U24580 ( .A(1'b0), .ZN(n35877) );
  INV_X1 U24582 ( .A(1'b0), .ZN(n35891) );
  INV_X1 U24584 ( .A(1'b0), .ZN(n35884) );
  INV_X1 U24586 ( .A(1'b0), .ZN(n35890) );
  INV_X1 U24588 ( .A(1'b0), .ZN(n35889) );
  INV_X1 U24590 ( .A(1'b0), .ZN(n35888) );
  INV_X1 U24592 ( .A(1'b0), .ZN(n35887) );
  INV_X1 U24594 ( .A(1'b0), .ZN(n35896) );
  INV_X1 U24596 ( .A(1'b0), .ZN(n35895) );
  INV_X1 U24598 ( .A(1'b0), .ZN(n33926) );
  INV_X1 U24600 ( .A(1'b0), .ZN(n35894) );
  INV_X1 U24602 ( .A(1'b0), .ZN(n35893) );
  INV_X1 U24604 ( .A(1'b0), .ZN(n33930) );
  INV_X1 U24606 ( .A(1'b0), .ZN(n35892) );
  INV_X1 U24608 ( .A(1'b0), .ZN(n35905) );
  INV_X1 U24610 ( .A(1'b0), .ZN(n35904) );
  INV_X1 U24612 ( .A(1'b0), .ZN(n35903) );
  INV_X1 U24614 ( .A(1'b0), .ZN(n35902) );
  INV_X1 U24616 ( .A(1'b0), .ZN(n35901) );
  INV_X1 U24618 ( .A(1'b0), .ZN(n35900) );
  INV_X1 U24620 ( .A(1'b0), .ZN(n35899) );
  INV_X1 U24622 ( .A(1'b0), .ZN(n35898) );
  INV_X1 U24624 ( .A(1'b0), .ZN(n35913) );
  INV_X1 U24626 ( .A(1'b0), .ZN(n35912) );
  INV_X1 U24628 ( .A(1'b0), .ZN(n35911) );
  INV_X1 U24630 ( .A(1'b0), .ZN(n35910) );
  INV_X1 U24632 ( .A(1'b0), .ZN(n35909) );
  INV_X1 U24634 ( .A(1'b0), .ZN(n35908) );
  INV_X1 U24636 ( .A(1'b0), .ZN(n35907) );
  INV_X1 U24638 ( .A(1'b0), .ZN(n35906) );
  INV_X1 U24640 ( .A(1'b0), .ZN(n35921) );
  INV_X1 U24642 ( .A(1'b0), .ZN(n35920) );
  INV_X1 U24644 ( .A(1'b0), .ZN(n35919) );
  INV_X1 U24646 ( .A(1'b0), .ZN(n35918) );
  INV_X1 U24648 ( .A(1'b0), .ZN(n35917) );
  INV_X1 U24650 ( .A(1'b0), .ZN(n35916) );
  INV_X1 U24652 ( .A(1'b0), .ZN(n35915) );
  INV_X1 U24654 ( .A(1'b0), .ZN(n35914) );
  INV_X1 U24656 ( .A(1'b0), .ZN(n35929) );
  INV_X1 U24658 ( .A(1'b0), .ZN(n35928) );
  INV_X1 U24660 ( .A(1'b0), .ZN(n35927) );
  INV_X1 U24662 ( .A(1'b0), .ZN(n35926) );
  INV_X1 U24664 ( .A(1'b0), .ZN(n35925) );
  INV_X1 U24666 ( .A(1'b0), .ZN(n35924) );
  INV_X1 U24668 ( .A(1'b0), .ZN(n35923) );
  INV_X1 U24670 ( .A(1'b0), .ZN(n35922) );
  INV_X1 U24672 ( .A(1'b0), .ZN(n35937) );
  INV_X1 U24674 ( .A(1'b0), .ZN(n35936) );
  INV_X1 U24676 ( .A(1'b0), .ZN(n35935) );
  INV_X1 U24678 ( .A(1'b0), .ZN(n35934) );
  INV_X1 U24680 ( .A(1'b0), .ZN(n35933) );
  INV_X1 U24682 ( .A(1'b0), .ZN(n35932) );
  INV_X1 U24684 ( .A(1'b0), .ZN(n35931) );
  INV_X1 U24686 ( .A(1'b0), .ZN(n35930) );
  INV_X1 U24688 ( .A(1'b0), .ZN(n35945) );
  INV_X1 U24690 ( .A(1'b0), .ZN(n35944) );
  INV_X1 U24692 ( .A(1'b0), .ZN(n35943) );
  INV_X1 U24694 ( .A(1'b0), .ZN(n35942) );
  INV_X1 U24696 ( .A(1'b0), .ZN(n35941) );
  INV_X1 U24698 ( .A(1'b0), .ZN(n35940) );
  INV_X1 U24700 ( .A(1'b0), .ZN(n35939) );
  INV_X1 U24702 ( .A(1'b0), .ZN(n35938) );
  INV_X1 U24704 ( .A(1'b0), .ZN(n35953) );
  INV_X1 U24706 ( .A(1'b0), .ZN(n35952) );
  INV_X1 U24708 ( .A(1'b0), .ZN(n35951) );
  INV_X1 U24710 ( .A(1'b0), .ZN(n35950) );
  INV_X1 U24712 ( .A(1'b0), .ZN(n35949) );
  INV_X1 U24714 ( .A(1'b0), .ZN(n35948) );
  INV_X1 U24716 ( .A(1'b0), .ZN(n35947) );
  INV_X1 U24718 ( .A(1'b0), .ZN(n35946) );
  INV_X1 U24720 ( .A(1'b0), .ZN(n35961) );
  INV_X1 U24722 ( .A(1'b0), .ZN(n35960) );
  INV_X1 U24724 ( .A(1'b0), .ZN(n35959) );
  INV_X1 U24726 ( .A(1'b0), .ZN(n35958) );
  INV_X1 U24728 ( .A(1'b0), .ZN(n35957) );
  INV_X1 U24730 ( .A(1'b0), .ZN(n35956) );
  INV_X1 U24732 ( .A(1'b0), .ZN(n35955) );
  INV_X1 U24734 ( .A(1'b0), .ZN(n35954) );
  INV_X1 U24736 ( .A(1'b0), .ZN(n35969) );
  INV_X1 U24738 ( .A(1'b0), .ZN(n35968) );
  INV_X1 U24740 ( .A(1'b0), .ZN(n35967) );
  INV_X1 U24742 ( .A(1'b0), .ZN(n35966) );
  INV_X1 U24744 ( .A(1'b0), .ZN(n35965) );
  INV_X1 U24746 ( .A(1'b0), .ZN(n35964) );
  INV_X1 U24748 ( .A(1'b0), .ZN(n35963) );
  INV_X1 U24750 ( .A(1'b0), .ZN(n35962) );
  INV_X1 U24752 ( .A(1'b0), .ZN(n35977) );
  INV_X1 U24754 ( .A(1'b0), .ZN(n35976) );
  INV_X1 U24756 ( .A(1'b0), .ZN(n35975) );
  INV_X1 U24758 ( .A(1'b0), .ZN(n35974) );
  INV_X1 U24760 ( .A(1'b0), .ZN(n35973) );
  INV_X1 U24762 ( .A(1'b0), .ZN(n35972) );
  INV_X1 U24764 ( .A(1'b0), .ZN(n35971) );
  INV_X1 U24766 ( .A(1'b0), .ZN(n35970) );
  INV_X1 U24768 ( .A(1'b0), .ZN(n35985) );
  INV_X1 U24770 ( .A(1'b0), .ZN(n35984) );
  INV_X1 U24772 ( .A(1'b0), .ZN(n35983) );
  INV_X1 U24774 ( .A(1'b0), .ZN(n35982) );
  INV_X1 U24776 ( .A(1'b0), .ZN(n35981) );
  INV_X1 U24778 ( .A(1'b0), .ZN(n35980) );
  INV_X1 U24780 ( .A(1'b0), .ZN(n35979) );
  INV_X1 U24782 ( .A(1'b0), .ZN(n35978) );
  INV_X1 U24784 ( .A(1'b0), .ZN(n35993) );
  INV_X1 U24786 ( .A(1'b0), .ZN(n35992) );
  INV_X1 U24788 ( .A(1'b0), .ZN(n35991) );
  INV_X1 U24790 ( .A(1'b0), .ZN(n35990) );
  INV_X1 U24792 ( .A(1'b0), .ZN(n35989) );
  INV_X1 U24794 ( .A(1'b0), .ZN(n35988) );
  INV_X1 U24796 ( .A(1'b0), .ZN(n35987) );
  INV_X1 U24798 ( .A(1'b0), .ZN(n35986) );
  INV_X1 U24800 ( .A(1'b0), .ZN(n36001) );
  INV_X1 U24802 ( .A(1'b0), .ZN(n36000) );
  INV_X1 U24804 ( .A(1'b0), .ZN(n35999) );
  INV_X1 U24806 ( .A(1'b0), .ZN(n35998) );
  INV_X1 U24808 ( .A(1'b0), .ZN(n35997) );
  INV_X1 U24810 ( .A(1'b0), .ZN(n35996) );
  INV_X1 U24812 ( .A(1'b0), .ZN(n35995) );
  INV_X1 U24814 ( .A(1'b0), .ZN(n35994) );
  INV_X1 U24816 ( .A(1'b0), .ZN(n36009) );
  INV_X1 U24818 ( .A(1'b0), .ZN(n36008) );
  INV_X1 U24820 ( .A(1'b0), .ZN(n36007) );
  INV_X1 U24822 ( .A(1'b0), .ZN(n36006) );
  INV_X1 U24824 ( .A(1'b0), .ZN(n36005) );
  INV_X1 U24826 ( .A(1'b0), .ZN(n36004) );
  INV_X1 U24828 ( .A(1'b0), .ZN(n36003) );
  INV_X1 U24830 ( .A(1'b0), .ZN(n36002) );
  INV_X1 U24832 ( .A(1'b0), .ZN(n36017) );
  INV_X1 U24834 ( .A(1'b0), .ZN(n36016) );
  INV_X1 U24836 ( .A(1'b0), .ZN(n36015) );
  INV_X1 U24838 ( .A(1'b0), .ZN(n36014) );
  INV_X1 U24840 ( .A(1'b0), .ZN(n36013) );
  INV_X1 U24842 ( .A(1'b0), .ZN(n36012) );
  INV_X1 U24844 ( .A(1'b0), .ZN(n36011) );
  INV_X1 U24846 ( .A(1'b0), .ZN(n36010) );
  INV_X1 U24848 ( .A(1'b0), .ZN(n36025) );
  INV_X1 U24850 ( .A(1'b0), .ZN(n36024) );
  INV_X1 U24852 ( .A(1'b0), .ZN(n36023) );
  INV_X1 U24854 ( .A(1'b0), .ZN(n36022) );
  INV_X1 U24856 ( .A(1'b0), .ZN(n36021) );
  INV_X1 U24858 ( .A(1'b0), .ZN(n36020) );
  INV_X1 U24860 ( .A(1'b0), .ZN(n36019) );
  INV_X1 U24862 ( .A(1'b0), .ZN(n36018) );
  INV_X1 U24864 ( .A(1'b0), .ZN(n36033) );
  INV_X1 U24866 ( .A(1'b0), .ZN(n36032) );
  INV_X1 U24868 ( .A(1'b0), .ZN(n36031) );
  INV_X1 U24870 ( .A(1'b0), .ZN(n36030) );
  INV_X1 U24872 ( .A(1'b0), .ZN(n36029) );
  INV_X1 U24874 ( .A(1'b0), .ZN(n36028) );
  INV_X1 U24876 ( .A(1'b0), .ZN(n36027) );
  INV_X1 U24878 ( .A(1'b0), .ZN(n36026) );
  INV_X1 U24880 ( .A(1'b0), .ZN(n36041) );
  INV_X1 U24882 ( .A(1'b0), .ZN(n36040) );
  INV_X1 U24884 ( .A(1'b0), .ZN(n36039) );
  INV_X1 U24886 ( .A(1'b0), .ZN(n36038) );
  INV_X1 U24888 ( .A(1'b0), .ZN(n36037) );
  INV_X1 U24890 ( .A(1'b0), .ZN(n36036) );
  INV_X1 U24892 ( .A(1'b0), .ZN(n36035) );
  INV_X1 U24894 ( .A(1'b0), .ZN(n36034) );
  INV_X1 U24896 ( .A(1'b0), .ZN(n36049) );
  INV_X1 U24898 ( .A(1'b0), .ZN(n36048) );
  INV_X1 U24900 ( .A(1'b0), .ZN(n36047) );
  INV_X1 U24902 ( .A(1'b0), .ZN(n36046) );
  INV_X1 U24904 ( .A(1'b0), .ZN(n36045) );
  INV_X1 U24906 ( .A(1'b0), .ZN(n36044) );
  INV_X1 U24908 ( .A(1'b0), .ZN(n36043) );
  INV_X1 U24910 ( .A(1'b0), .ZN(n36042) );
  INV_X1 U24912 ( .A(1'b0), .ZN(n36057) );
  INV_X1 U24914 ( .A(1'b0), .ZN(n36056) );
  INV_X1 U24916 ( .A(1'b0), .ZN(n36055) );
  INV_X1 U24918 ( .A(1'b0), .ZN(n36054) );
  INV_X1 U24920 ( .A(1'b0), .ZN(n36053) );
  INV_X1 U24922 ( .A(1'b0), .ZN(n36052) );
  INV_X1 U24924 ( .A(1'b0), .ZN(n36051) );
  INV_X1 U24926 ( .A(1'b0), .ZN(n36050) );
  INV_X1 U24928 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1753) );
  INV_X1 U24930 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1752) );
  INV_X1 U24932 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1751) );
  INV_X1 U24934 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1750) );
  INV_X1 U24936 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1749) );
  INV_X1 U24938 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1747) );
  INV_X1 U24940 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1746) );
  INV_X1 U24942 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1745) );
  INV_X1 U24944 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1743) );
  INV_X1 U24946 ( .A(1'b0), .ZN(p_wishbone_tx_fifo_n1742) );
  INV_X1 U24948 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1708) );
  INV_X1 U24950 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1707) );
  INV_X1 U24952 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1706) );
  INV_X1 U24954 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1705) );
  INV_X1 U24956 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1704) );
  INV_X1 U24958 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1703) );
  INV_X1 U24960 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1702) );
  INV_X1 U24962 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1701) );
  INV_X1 U24964 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1700) );
  INV_X1 U24966 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1699) );
  INV_X1 U24968 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1698) );
  INV_X1 U24970 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1697) );
  INV_X1 U24972 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1696) );
  INV_X1 U24974 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1695) );
  INV_X1 U24976 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1694) );
  INV_X1 U24978 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1693) );
  INV_X1 U24980 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1692) );
  INV_X1 U24982 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1691) );
  INV_X1 U24984 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1690) );
  INV_X1 U24986 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1689) );
  INV_X1 U24988 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1688) );
  INV_X1 U24990 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1687) );
  INV_X1 U24992 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1686) );
  INV_X1 U24994 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1685) );
  INV_X1 U24996 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1684) );
  INV_X1 U24998 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1683) );
  INV_X1 U25000 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1682) );
  INV_X1 U25002 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1681) );
  INV_X1 U25004 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1680) );
  INV_X1 U25006 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1679) );
  INV_X1 U25008 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1678) );
  INV_X1 U25010 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1677) );
  INV_X1 U25012 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1676) );
  INV_X1 U25014 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1675) );
  INV_X1 U25016 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1674) );
  INV_X1 U25018 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1673) );
  INV_X1 U25020 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1672) );
  INV_X1 U25022 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1671) );
  INV_X1 U25024 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1670) );
  INV_X1 U25026 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1669) );
  INV_X1 U25028 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1668) );
  INV_X1 U25030 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1667) );
  INV_X1 U25032 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1666) );
  INV_X1 U25034 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1665) );
  INV_X1 U25036 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1664) );
  INV_X1 U25038 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1663) );
  INV_X1 U25040 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1662) );
  INV_X1 U25042 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1661) );
  INV_X1 U25044 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1660) );
  INV_X1 U25046 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1659) );
  INV_X1 U25048 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1658) );
  INV_X1 U25050 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1657) );
  INV_X1 U25052 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1656) );
  INV_X1 U25054 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1655) );
  INV_X1 U25056 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1654) );
  INV_X1 U25058 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1653) );
  INV_X1 U25060 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1652) );
  INV_X1 U25062 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1651) );
  INV_X1 U25064 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1650) );
  INV_X1 U25066 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1649) );
  INV_X1 U25068 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1648) );
  INV_X1 U25070 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1647) );
  INV_X1 U25072 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1646) );
  INV_X1 U25074 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1645) );
  INV_X1 U25076 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1644) );
  INV_X1 U25078 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1643) );
  INV_X1 U25080 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1642) );
  INV_X1 U25082 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1641) );
  INV_X1 U25084 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1640) );
  INV_X1 U25086 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1639) );
  INV_X1 U25088 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1638) );
  INV_X1 U25090 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1637) );
  INV_X1 U25092 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1636) );
  INV_X1 U25094 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1635) );
  INV_X1 U25096 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1634) );
  INV_X1 U25098 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1633) );
  INV_X1 U25100 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1632) );
  INV_X1 U25102 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1631) );
  INV_X1 U25104 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1630) );
  INV_X1 U25106 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1629) );
  INV_X1 U25108 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1628) );
  INV_X1 U25110 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1627) );
  INV_X1 U25112 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1626) );
  INV_X1 U25114 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1625) );
  INV_X1 U25116 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1624) );
  INV_X1 U25118 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1623) );
  INV_X1 U25120 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1622) );
  INV_X1 U25122 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1621) );
  INV_X1 U25124 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1620) );
  INV_X1 U25126 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1619) );
  INV_X1 U25128 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1618) );
  INV_X1 U25130 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1617) );
  INV_X1 U25132 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1616) );
  INV_X1 U25134 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1615) );
  INV_X1 U25136 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1614) );
  INV_X1 U25138 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1613) );
  INV_X1 U25140 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1612) );
  INV_X1 U25142 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1611) );
  INV_X1 U25144 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1610) );
  INV_X1 U25146 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1609) );
  INV_X1 U25148 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1608) );
  INV_X1 U25150 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1607) );
  INV_X1 U25152 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1606) );
  INV_X1 U25154 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1605) );
  INV_X1 U25156 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1604) );
  INV_X1 U25158 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1603) );
  INV_X1 U25160 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1602) );
  INV_X1 U25162 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1601) );
  INV_X1 U25164 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1600) );
  INV_X1 U25166 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1599) );
  INV_X1 U25168 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1598) );
  INV_X1 U25170 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1597) );
  INV_X1 U25172 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1596) );
  INV_X1 U25174 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1595) );
  INV_X1 U25176 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1594) );
  INV_X1 U25178 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1593) );
  INV_X1 U25180 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1592) );
  INV_X1 U25182 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1591) );
  INV_X1 U25184 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1590) );
  INV_X1 U25186 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1589) );
  INV_X1 U25188 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1588) );
  INV_X1 U25190 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1587) );
  INV_X1 U25192 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1586) );
  INV_X1 U25194 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1585) );
  INV_X1 U25196 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1584) );
  INV_X1 U25198 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1583) );
  INV_X1 U25200 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1582) );
  INV_X1 U25202 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1581) );
  INV_X1 U25204 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1580) );
  INV_X1 U25206 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1579) );
  INV_X1 U25208 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1578) );
  INV_X1 U25210 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1577) );
  INV_X1 U25212 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1576) );
  INV_X1 U25214 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1575) );
  INV_X1 U25216 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1574) );
  INV_X1 U25218 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1573) );
  INV_X1 U25220 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1572) );
  INV_X1 U25222 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1571) );
  INV_X1 U25224 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1570) );
  INV_X1 U25226 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1569) );
  INV_X1 U25228 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1568) );
  INV_X1 U25230 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1567) );
  INV_X1 U25232 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1566) );
  INV_X1 U25234 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1565) );
  INV_X1 U25236 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1564) );
  INV_X1 U25238 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1563) );
  INV_X1 U25240 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1562) );
  INV_X1 U25242 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1561) );
  INV_X1 U25244 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1560) );
  INV_X1 U25246 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1559) );
  INV_X1 U25248 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1558) );
  INV_X1 U25250 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1557) );
  INV_X1 U25252 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1556) );
  INV_X1 U25254 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1555) );
  INV_X1 U25256 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1554) );
  INV_X1 U25258 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1553) );
  INV_X1 U25260 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1552) );
  INV_X1 U25262 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1551) );
  INV_X1 U25264 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1550) );
  INV_X1 U25266 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1549) );
  INV_X1 U25268 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1548) );
  INV_X1 U25270 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1547) );
  INV_X1 U25272 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1546) );
  INV_X1 U25274 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1545) );
  INV_X1 U25276 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1544) );
  INV_X1 U25278 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1543) );
  INV_X1 U25280 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1542) );
  INV_X1 U25282 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1541) );
  INV_X1 U25284 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1540) );
  INV_X1 U25286 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1539) );
  INV_X1 U25288 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1538) );
  INV_X1 U25290 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1537) );
  INV_X1 U25292 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1536) );
  INV_X1 U25294 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1535) );
  INV_X1 U25296 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1534) );
  INV_X1 U25298 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1533) );
  INV_X1 U25300 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1532) );
  INV_X1 U25302 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1531) );
  INV_X1 U25304 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1530) );
  INV_X1 U25306 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1529) );
  INV_X1 U25308 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1528) );
  INV_X1 U25310 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1527) );
  INV_X1 U25312 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1526) );
  INV_X1 U25314 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1525) );
  INV_X1 U25316 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1524) );
  INV_X1 U25318 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1523) );
  INV_X1 U25320 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1522) );
  INV_X1 U25322 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1521) );
  INV_X1 U25324 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1520) );
  INV_X1 U25326 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1519) );
  INV_X1 U25328 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1518) );
  INV_X1 U25330 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1517) );
  INV_X1 U25332 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1516) );
  INV_X1 U25334 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1515) );
  INV_X1 U25336 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1514) );
  INV_X1 U25338 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1513) );
  INV_X1 U25340 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1512) );
  INV_X1 U25342 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1511) );
  INV_X1 U25344 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1510) );
  INV_X1 U25346 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1509) );
  INV_X1 U25348 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1508) );
  INV_X1 U25350 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1507) );
  INV_X1 U25352 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1506) );
  INV_X1 U25354 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1505) );
  INV_X1 U25356 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1504) );
  INV_X1 U25358 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1503) );
  INV_X1 U25360 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1502) );
  INV_X1 U25362 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1501) );
  INV_X1 U25364 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1500) );
  INV_X1 U25366 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1499) );
  INV_X1 U25368 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1498) );
  INV_X1 U25370 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1497) );
  INV_X1 U25372 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1496) );
  INV_X1 U25374 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1495) );
  INV_X1 U25376 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1494) );
  INV_X1 U25378 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1493) );
  INV_X1 U25380 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1492) );
  INV_X1 U25382 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1491) );
  INV_X1 U25384 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1490) );
  INV_X1 U25386 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1489) );
  INV_X1 U25388 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1488) );
  INV_X1 U25390 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1487) );
  INV_X1 U25392 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1486) );
  INV_X1 U25394 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1485) );
  INV_X1 U25396 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1484) );
  INV_X1 U25398 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1483) );
  INV_X1 U25400 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1482) );
  INV_X1 U25402 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1481) );
  INV_X1 U25404 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1480) );
  INV_X1 U25406 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1479) );
  INV_X1 U25408 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1478) );
  INV_X1 U25410 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1477) );
  INV_X1 U25412 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1476) );
  INV_X1 U25414 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1475) );
  INV_X1 U25416 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1474) );
  INV_X1 U25418 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1473) );
  INV_X1 U25420 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1472) );
  INV_X1 U25422 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1471) );
  INV_X1 U25424 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1470) );
  INV_X1 U25426 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1469) );
  INV_X1 U25428 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1468) );
  INV_X1 U25430 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1467) );
  INV_X1 U25432 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1466) );
  INV_X1 U25434 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1465) );
  INV_X1 U25436 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1464) );
  INV_X1 U25438 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1463) );
  INV_X1 U25440 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1462) );
  INV_X1 U25442 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1461) );
  INV_X1 U25444 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1460) );
  INV_X1 U25446 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1459) );
  INV_X1 U25448 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1458) );
  INV_X1 U25450 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1457) );
  INV_X1 U25452 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1456) );
  INV_X1 U25454 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1455) );
  INV_X1 U25456 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1454) );
  INV_X1 U25458 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1453) );
  INV_X1 U25460 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1452) );
  INV_X1 U25462 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1451) );
  INV_X1 U25464 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1450) );
  INV_X1 U25466 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1449) );
  INV_X1 U25468 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1448) );
  INV_X1 U25470 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1447) );
  INV_X1 U25472 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1446) );
  INV_X1 U25474 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1445) );
  INV_X1 U25476 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1444) );
  INV_X1 U25478 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1443) );
  INV_X1 U25480 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1442) );
  INV_X1 U25482 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1441) );
  INV_X1 U25484 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1440) );
  INV_X1 U25486 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1439) );
  INV_X1 U25488 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1438) );
  INV_X1 U25490 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1437) );
  INV_X1 U25492 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1436) );
  INV_X1 U25494 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1435) );
  INV_X1 U25496 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1434) );
  INV_X1 U25498 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1433) );
  INV_X1 U25500 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1432) );
  INV_X1 U25502 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1431) );
  INV_X1 U25504 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1430) );
  INV_X1 U25506 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1429) );
  INV_X1 U25508 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1428) );
  INV_X1 U25510 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1427) );
  INV_X1 U25512 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1426) );
  INV_X1 U25514 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1425) );
  INV_X1 U25516 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1424) );
  INV_X1 U25518 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1423) );
  INV_X1 U25520 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1422) );
  INV_X1 U25522 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1421) );
  INV_X1 U25524 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1420) );
  INV_X1 U25526 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1419) );
  INV_X1 U25528 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1418) );
  INV_X1 U25530 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1417) );
  INV_X1 U25532 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1416) );
  INV_X1 U25534 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1415) );
  INV_X1 U25536 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1414) );
  INV_X1 U25538 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1413) );
  INV_X1 U25540 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1412) );
  INV_X1 U25542 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1411) );
  INV_X1 U25544 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1410) );
  INV_X1 U25546 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1409) );
  INV_X1 U25548 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1408) );
  INV_X1 U25550 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1407) );
  INV_X1 U25552 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1406) );
  INV_X1 U25554 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1405) );
  INV_X1 U25556 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1404) );
  INV_X1 U25558 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1403) );
  INV_X1 U25560 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1402) );
  INV_X1 U25562 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1401) );
  INV_X1 U25564 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1400) );
  INV_X1 U25566 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1399) );
  INV_X1 U25568 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1398) );
  INV_X1 U25570 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1397) );
  INV_X1 U25572 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1396) );
  INV_X1 U25574 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1395) );
  INV_X1 U25576 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1394) );
  INV_X1 U25578 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1393) );
  INV_X1 U25580 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1392) );
  INV_X1 U25582 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1391) );
  INV_X1 U25584 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1390) );
  INV_X1 U25586 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1389) );
  INV_X1 U25588 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1388) );
  INV_X1 U25590 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1387) );
  INV_X1 U25592 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1386) );
  INV_X1 U25594 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1385) );
  INV_X1 U25596 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1384) );
  INV_X1 U25598 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1383) );
  INV_X1 U25600 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1382) );
  INV_X1 U25602 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1381) );
  INV_X1 U25604 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1380) );
  INV_X1 U25606 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1379) );
  INV_X1 U25608 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1378) );
  INV_X1 U25610 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1377) );
  INV_X1 U25612 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1376) );
  INV_X1 U25614 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1375) );
  INV_X1 U25616 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1374) );
  INV_X1 U25618 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1373) );
  INV_X1 U25620 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1372) );
  INV_X1 U25622 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1371) );
  INV_X1 U25624 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1370) );
  INV_X1 U25626 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1369) );
  INV_X1 U25628 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1368) );
  INV_X1 U25630 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1367) );
  INV_X1 U25632 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1366) );
  INV_X1 U25634 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1365) );
  INV_X1 U25636 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1364) );
  INV_X1 U25638 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1363) );
  INV_X1 U25640 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1362) );
  INV_X1 U25642 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1361) );
  INV_X1 U25644 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1360) );
  INV_X1 U25646 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1359) );
  INV_X1 U25648 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1358) );
  INV_X1 U25650 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1357) );
  INV_X1 U25652 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1356) );
  INV_X1 U25654 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1355) );
  INV_X1 U25656 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1354) );
  INV_X1 U25658 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1353) );
  INV_X1 U25660 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1352) );
  INV_X1 U25662 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1351) );
  INV_X1 U25664 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1350) );
  INV_X1 U25666 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1349) );
  INV_X1 U25668 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1348) );
  INV_X1 U25670 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1347) );
  INV_X1 U25672 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1346) );
  INV_X1 U25674 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1345) );
  INV_X1 U25676 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1344) );
  INV_X1 U25678 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1343) );
  INV_X1 U25680 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1342) );
  INV_X1 U25682 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1341) );
  INV_X1 U25684 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1340) );
  INV_X1 U25686 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1339) );
  INV_X1 U25688 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1338) );
  INV_X1 U25690 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1337) );
  INV_X1 U25692 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1336) );
  INV_X1 U25694 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1335) );
  INV_X1 U25696 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1334) );
  INV_X1 U25698 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1333) );
  INV_X1 U25700 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1332) );
  INV_X1 U25702 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1331) );
  INV_X1 U25704 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1330) );
  INV_X1 U25706 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1329) );
  INV_X1 U25708 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1328) );
  INV_X1 U25710 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1327) );
  INV_X1 U25712 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1326) );
  INV_X1 U25714 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1325) );
  INV_X1 U25716 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1324) );
  INV_X1 U25718 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1323) );
  INV_X1 U25720 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1322) );
  INV_X1 U25722 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1321) );
  INV_X1 U25724 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1320) );
  INV_X1 U25726 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1319) );
  INV_X1 U25728 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1318) );
  INV_X1 U25730 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1317) );
  INV_X1 U25732 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1316) );
  INV_X1 U25734 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1315) );
  INV_X1 U25736 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1314) );
  INV_X1 U25738 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1313) );
  INV_X1 U25740 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1312) );
  INV_X1 U25742 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1311) );
  INV_X1 U25744 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1310) );
  INV_X1 U25746 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1309) );
  INV_X1 U25748 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1308) );
  INV_X1 U25750 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1307) );
  INV_X1 U25752 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1306) );
  INV_X1 U25754 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1305) );
  INV_X1 U25756 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1304) );
  INV_X1 U25758 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1303) );
  INV_X1 U25760 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1302) );
  INV_X1 U25762 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1301) );
  INV_X1 U25764 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1300) );
  INV_X1 U25766 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1299) );
  INV_X1 U25768 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1298) );
  INV_X1 U25770 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1297) );
  INV_X1 U25772 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1296) );
  INV_X1 U25774 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1295) );
  INV_X1 U25776 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1294) );
  INV_X1 U25778 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1293) );
  INV_X1 U25780 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1292) );
  INV_X1 U25782 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1291) );
  INV_X1 U25784 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1290) );
  INV_X1 U25786 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1289) );
  INV_X1 U25788 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1288) );
  INV_X1 U25790 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1287) );
  INV_X1 U25792 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1286) );
  INV_X1 U25794 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1285) );
  INV_X1 U25796 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1284) );
  INV_X1 U25798 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1283) );
  INV_X1 U25800 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1282) );
  INV_X1 U25802 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1281) );
  INV_X1 U25804 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1280) );
  INV_X1 U25806 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1279) );
  INV_X1 U25808 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1278) );
  INV_X1 U25810 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1277) );
  INV_X1 U25812 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1276) );
  INV_X1 U25814 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1275) );
  INV_X1 U25816 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1274) );
  INV_X1 U25818 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1273) );
  INV_X1 U25820 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1272) );
  INV_X1 U25822 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1271) );
  INV_X1 U25824 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1270) );
  INV_X1 U25826 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1269) );
  INV_X1 U25828 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1268) );
  INV_X1 U25830 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1267) );
  INV_X1 U25832 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1266) );
  INV_X1 U25834 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1265) );
  INV_X1 U25836 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1264) );
  INV_X1 U25838 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1263) );
  INV_X1 U25840 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1262) );
  INV_X1 U25842 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1261) );
  INV_X1 U25844 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1260) );
  INV_X1 U25846 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1259) );
  INV_X1 U25848 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1258) );
  INV_X1 U25850 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1257) );
  INV_X1 U25852 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1256) );
  INV_X1 U25854 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1255) );
  INV_X1 U25856 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1254) );
  INV_X1 U25858 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1253) );
  INV_X1 U25860 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1252) );
  INV_X1 U25862 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1251) );
  INV_X1 U25864 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1250) );
  INV_X1 U25866 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1249) );
  INV_X1 U25868 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1248) );
  INV_X1 U25870 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1247) );
  INV_X1 U25872 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1246) );
  INV_X1 U25874 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1245) );
  INV_X1 U25876 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1244) );
  INV_X1 U25878 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1243) );
  INV_X1 U25880 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1242) );
  INV_X1 U25882 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1241) );
  INV_X1 U25884 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1240) );
  INV_X1 U25886 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1239) );
  INV_X1 U25888 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1238) );
  INV_X1 U25890 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1237) );
  INV_X1 U25892 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1236) );
  INV_X1 U25894 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1235) );
  INV_X1 U25896 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1234) );
  INV_X1 U25898 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1233) );
  INV_X1 U25900 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1232) );
  INV_X1 U25902 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1231) );
  INV_X1 U25904 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1230) );
  INV_X1 U25906 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_n1229) );
  INV_X1 U25908 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N654) );
  INV_X1 U25910 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N653) );
  INV_X1 U25912 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N652) );
  INV_X1 U25914 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N651) );
  INV_X1 U25916 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N650) );
  INV_X1 U25918 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N649) );
  INV_X1 U25920 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N648) );
  INV_X1 U25922 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N647) );
  INV_X1 U25924 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N646) );
  INV_X1 U25926 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N645) );
  INV_X1 U25928 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N644) );
  INV_X1 U25930 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N643) );
  INV_X1 U25932 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N642) );
  INV_X1 U25934 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N641) );
  INV_X1 U25936 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N640) );
  INV_X1 U25938 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N639) );
  INV_X1 U25940 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N638) );
  INV_X1 U25942 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N637) );
  INV_X1 U25944 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N636) );
  INV_X1 U25946 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N635) );
  INV_X1 U25948 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N634) );
  INV_X1 U25950 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N633) );
  INV_X1 U25952 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N632) );
  INV_X1 U25954 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N631) );
  INV_X1 U25956 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N630) );
  INV_X1 U25958 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N629) );
  INV_X1 U25960 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N628) );
  INV_X1 U25962 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N627) );
  INV_X1 U25964 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N626) );
  INV_X1 U25966 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N625) );
  INV_X1 U25968 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N624) );
  INV_X1 U25970 ( .A(1'b1), .ZN(p_wishbone_tx_fifo_N623) );
  INV_X1 U25972 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25360) );
  INV_X1 U25974 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25358) );
  INV_X1 U25976 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25355) );
  INV_X1 U25978 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25353) );
  INV_X1 U25980 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25311) );
  INV_X1 U25982 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25309) );
  INV_X1 U25984 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25308) );
  INV_X1 U25986 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25306) );
  INV_X1 U25988 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25264) );
  INV_X1 U25990 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25262) );
  INV_X1 U25992 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25259) );
  INV_X1 U25994 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25257) );
  INV_X1 U25996 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25208) );
  INV_X1 U25998 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25206) );
  INV_X1 U26000 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25203) );
  INV_X1 U26002 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25201) );
  INV_X1 U26004 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25136) );
  INV_X1 U26006 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25134) );
  INV_X1 U26008 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25131) );
  INV_X1 U26010 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25129) );
  INV_X1 U26012 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n25000) );
  INV_X1 U26014 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24998) );
  INV_X1 U26016 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24995) );
  INV_X1 U26018 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24993) );
  INV_X1 U26020 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24992) );
  INV_X1 U26022 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24990) );
  INV_X1 U26024 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24987) );
  INV_X1 U26026 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24985) );
  INV_X1 U26028 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24968) );
  INV_X1 U26030 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24966) );
  INV_X1 U26032 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24963) );
  INV_X1 U26034 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24961) );
  INV_X1 U26036 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24920) );
  INV_X1 U26038 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24918) );
  INV_X1 U26040 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24915) );
  INV_X1 U26042 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24913) );
  INV_X1 U26044 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24896) );
  INV_X1 U26046 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24894) );
  INV_X1 U26048 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24891) );
  INV_X1 U26050 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24889) );
  INV_X1 U26052 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24832) );
  INV_X1 U26054 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24830) );
  INV_X1 U26056 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24827) );
  INV_X1 U26058 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24825) );
  INV_X1 U26060 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24824) );
  INV_X1 U26062 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24822) );
  INV_X1 U26064 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24819) );
  INV_X1 U26066 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24817) );
  INV_X1 U26068 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24808) );
  INV_X1 U26070 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24806) );
  INV_X1 U26072 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24803) );
  INV_X1 U26074 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24801) );
  INV_X1 U26076 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24768) );
  INV_X1 U26078 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24766) );
  INV_X1 U26080 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24763) );
  INV_X1 U26082 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24761) );
  INV_X1 U26084 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24704) );
  INV_X1 U26086 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24702) );
  INV_X1 U26088 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24699) );
  INV_X1 U26090 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24697) );
  INV_X1 U26092 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24680) );
  INV_X1 U26094 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24678) );
  INV_X1 U26096 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24675) );
  INV_X1 U26098 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24673) );
  INV_X1 U26100 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24608) );
  INV_X1 U26102 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24606) );
  INV_X1 U26104 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24603) );
  INV_X1 U26106 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24601) );
  INV_X1 U26108 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24584) );
  INV_X1 U26110 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24582) );
  INV_X1 U26112 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24579) );
  INV_X1 U26114 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24577) );
  INV_X1 U26116 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24528) );
  INV_X1 U26118 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24526) );
  INV_X1 U26120 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24523) );
  INV_X1 U26122 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24521) );
  INV_X1 U26124 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24520) );
  INV_X1 U26126 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24518) );
  INV_X1 U26128 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24515) );
  INV_X1 U26130 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24513) );
  INV_X1 U26132 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24368) );
  INV_X1 U26134 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24366) );
  INV_X1 U26136 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24363) );
  INV_X1 U26138 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24361) );
  INV_X1 U26140 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24351) );
  INV_X1 U26142 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24349) );
  INV_X1 U26144 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24348) );
  INV_X1 U26146 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24346) );
  INV_X1 U26148 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24295) );
  INV_X1 U26150 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24293) );
  INV_X1 U26152 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24292) );
  INV_X1 U26154 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24290) );
  INV_X1 U26156 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24264) );
  INV_X1 U26158 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24262) );
  INV_X1 U26160 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24259) );
  INV_X1 U26162 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24257) );
  INV_X1 U26164 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24199) );
  INV_X1 U26166 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24197) );
  INV_X1 U26168 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24196) );
  INV_X1 U26170 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24194) );
  INV_X1 U26172 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24184) );
  INV_X1 U26174 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24182) );
  INV_X1 U26176 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24179) );
  INV_X1 U26178 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24177) );
  INV_X1 U26180 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24176) );
  INV_X1 U26182 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24174) );
  INV_X1 U26184 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24171) );
  INV_X1 U26186 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24169) );
  INV_X1 U26188 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24168) );
  INV_X1 U26190 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24166) );
  INV_X1 U26192 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24163) );
  INV_X1 U26194 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24161) );
  INV_X1 U26196 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24136) );
  INV_X1 U26198 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24134) );
  INV_X1 U26200 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24131) );
  INV_X1 U26202 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24129) );
  INV_X1 U26204 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24119) );
  INV_X1 U26206 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24117) );
  INV_X1 U26208 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24116) );
  INV_X1 U26210 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24114) );
  INV_X1 U26212 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24103) );
  INV_X1 U26214 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24101) );
  INV_X1 U26216 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24100) );
  INV_X1 U26218 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24098) );
  INV_X1 U26220 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24088) );
  INV_X1 U26222 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24086) );
  INV_X1 U26224 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24083) );
  INV_X1 U26226 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24081) );
  INV_X1 U26228 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24079) );
  INV_X1 U26230 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24077) );
  INV_X1 U26232 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24076) );
  INV_X1 U26234 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24074) );
  INV_X1 U26236 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24071) );
  INV_X1 U26238 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24069) );
  INV_X1 U26240 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24068) );
  INV_X1 U26242 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24066) );
  INV_X1 U26244 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24063) );
  INV_X1 U26246 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24061) );
  INV_X1 U26248 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24060) );
  INV_X1 U26250 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24058) );
  INV_X1 U26252 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24056) );
  INV_X1 U26254 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24054) );
  INV_X1 U26256 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24051) );
  INV_X1 U26258 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24049) );
  INV_X1 U26260 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24024) );
  INV_X1 U26262 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24022) );
  INV_X1 U26264 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24019) );
  INV_X1 U26266 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24017) );
  INV_X1 U26268 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n24000) );
  INV_X1 U26270 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23998) );
  INV_X1 U26272 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23995) );
  INV_X1 U26274 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23993) );
  INV_X1 U26276 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23992) );
  INV_X1 U26278 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23990) );
  INV_X1 U26280 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23987) );
  INV_X1 U26282 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23985) );
  INV_X1 U26284 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23312) );
  INV_X1 U26286 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23310) );
  INV_X1 U26288 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23307) );
  INV_X1 U26290 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23305) );
  INV_X1 U26292 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23263) );
  INV_X1 U26294 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23261) );
  INV_X1 U26296 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23260) );
  INV_X1 U26298 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23258) );
  INV_X1 U26300 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23216) );
  INV_X1 U26302 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23214) );
  INV_X1 U26304 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23211) );
  INV_X1 U26306 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23209) );
  INV_X1 U26308 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23160) );
  INV_X1 U26310 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23158) );
  INV_X1 U26312 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23155) );
  INV_X1 U26314 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23153) );
  INV_X1 U26316 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23088) );
  INV_X1 U26318 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23086) );
  INV_X1 U26320 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23083) );
  INV_X1 U26322 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23081) );
  INV_X1 U26324 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23024) );
  INV_X1 U26326 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23022) );
  INV_X1 U26328 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23019) );
  INV_X1 U26330 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n23017) );
  INV_X1 U26332 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22976) );
  INV_X1 U26334 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22974) );
  INV_X1 U26336 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22971) );
  INV_X1 U26338 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22969) );
  INV_X1 U26340 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22952) );
  INV_X1 U26342 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22950) );
  INV_X1 U26344 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22947) );
  INV_X1 U26346 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22945) );
  INV_X1 U26348 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22888) );
  INV_X1 U26350 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22886) );
  INV_X1 U26352 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22883) );
  INV_X1 U26354 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22881) );
  INV_X1 U26356 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22880) );
  INV_X1 U26358 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22878) );
  INV_X1 U26360 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22875) );
  INV_X1 U26362 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22873) );
  INV_X1 U26364 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22864) );
  INV_X1 U26366 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22862) );
  INV_X1 U26368 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22859) );
  INV_X1 U26370 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22857) );
  INV_X1 U26372 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22824) );
  INV_X1 U26374 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22822) );
  INV_X1 U26376 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22819) );
  INV_X1 U26378 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22817) );
  INV_X1 U26380 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22760) );
  INV_X1 U26382 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22758) );
  INV_X1 U26384 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22755) );
  INV_X1 U26386 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22753) );
  INV_X1 U26388 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22736) );
  INV_X1 U26390 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22734) );
  INV_X1 U26392 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22731) );
  INV_X1 U26394 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22729) );
  INV_X1 U26396 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22664) );
  INV_X1 U26398 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22662) );
  INV_X1 U26400 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22659) );
  INV_X1 U26402 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22657) );
  INV_X1 U26404 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22640) );
  INV_X1 U26406 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22638) );
  INV_X1 U26408 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22635) );
  INV_X1 U26410 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22633) );
  INV_X1 U26412 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22584) );
  INV_X1 U26414 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22582) );
  INV_X1 U26416 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22579) );
  INV_X1 U26418 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22577) );
  INV_X1 U26420 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22576) );
  INV_X1 U26422 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22574) );
  INV_X1 U26424 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22571) );
  INV_X1 U26426 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22569) );
  INV_X1 U26428 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22440) );
  INV_X1 U26430 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22438) );
  INV_X1 U26432 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22435) );
  INV_X1 U26434 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22433) );
  INV_X1 U26436 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22432) );
  INV_X1 U26438 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22430) );
  INV_X1 U26440 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22427) );
  INV_X1 U26442 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22425) );
  INV_X1 U26444 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22328) );
  INV_X1 U26446 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22326) );
  INV_X1 U26448 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22323) );
  INV_X1 U26450 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22321) );
  INV_X1 U26452 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22312) );
  INV_X1 U26454 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22310) );
  INV_X1 U26456 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22307) );
  INV_X1 U26458 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22305) );
  INV_X1 U26460 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22264) );
  INV_X1 U26462 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22262) );
  INV_X1 U26464 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22259) );
  INV_X1 U26466 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22257) );
  INV_X1 U26468 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22232) );
  INV_X1 U26470 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22230) );
  INV_X1 U26472 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22227) );
  INV_X1 U26474 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22225) );
  INV_X1 U26476 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22208) );
  INV_X1 U26478 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22206) );
  INV_X1 U26480 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22203) );
  INV_X1 U26482 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22201) );
  INV_X1 U26484 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22168) );
  INV_X1 U26486 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22166) );
  INV_X1 U26488 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22163) );
  INV_X1 U26490 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22161) );
  INV_X1 U26492 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22151) );
  INV_X1 U26494 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22149) );
  INV_X1 U26496 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22148) );
  INV_X1 U26498 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22146) );
  INV_X1 U26500 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22144) );
  INV_X1 U26502 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22142) );
  INV_X1 U26504 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22139) );
  INV_X1 U26506 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22137) );
  INV_X1 U26508 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22136) );
  INV_X1 U26510 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22134) );
  INV_X1 U26512 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22131) );
  INV_X1 U26514 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22129) );
  INV_X1 U26516 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22112) );
  INV_X1 U26518 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22110) );
  INV_X1 U26520 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22107) );
  INV_X1 U26522 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22105) );
  INV_X1 U26524 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22104) );
  INV_X1 U26526 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22102) );
  INV_X1 U26528 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22099) );
  INV_X1 U26530 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22097) );
  INV_X1 U26532 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22096) );
  INV_X1 U26534 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22094) );
  INV_X1 U26536 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22091) );
  INV_X1 U26538 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22089) );
  INV_X1 U26540 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22080) );
  INV_X1 U26542 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22078) );
  INV_X1 U26544 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22075) );
  INV_X1 U26546 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22073) );
  INV_X1 U26548 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22064) );
  INV_X1 U26550 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22062) );
  INV_X1 U26552 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22059) );
  INV_X1 U26554 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22057) );
  INV_X1 U26556 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22048) );
  INV_X1 U26558 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22046) );
  INV_X1 U26560 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22043) );
  INV_X1 U26562 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22041) );
  INV_X1 U26564 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22040) );
  INV_X1 U26566 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22038) );
  INV_X1 U26568 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22035) );
  INV_X1 U26570 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22033) );
  INV_X1 U26572 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22023) );
  INV_X1 U26574 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22021) );
  INV_X1 U26576 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22020) );
  INV_X1 U26578 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22018) );
  INV_X1 U26580 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22015) );
  INV_X1 U26582 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22013) );
  INV_X1 U26584 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22012) );
  INV_X1 U26586 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n22010) );
  INV_X1 U26588 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21984) );
  INV_X1 U26590 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21982) );
  INV_X1 U26592 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21979) );
  INV_X1 U26594 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21977) );
  INV_X1 U26596 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21264) );
  INV_X1 U26598 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21262) );
  INV_X1 U26600 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21259) );
  INV_X1 U26602 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21257) );
  INV_X1 U26604 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21215) );
  INV_X1 U26606 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21213) );
  INV_X1 U26608 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21212) );
  INV_X1 U26610 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21210) );
  INV_X1 U26612 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21168) );
  INV_X1 U26614 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21166) );
  INV_X1 U26616 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21163) );
  INV_X1 U26618 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21161) );
  INV_X1 U26620 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21112) );
  INV_X1 U26622 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21110) );
  INV_X1 U26624 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21107) );
  INV_X1 U26626 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21105) );
  INV_X1 U26628 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21040) );
  INV_X1 U26630 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21038) );
  INV_X1 U26632 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21035) );
  INV_X1 U26634 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n21033) );
  INV_X1 U26636 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20976) );
  INV_X1 U26638 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20974) );
  INV_X1 U26640 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20971) );
  INV_X1 U26642 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20969) );
  INV_X1 U26644 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20928) );
  INV_X1 U26646 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20926) );
  INV_X1 U26648 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20923) );
  INV_X1 U26650 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20921) );
  INV_X1 U26652 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20904) );
  INV_X1 U26654 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20902) );
  INV_X1 U26656 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20899) );
  INV_X1 U26658 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20897) );
  INV_X1 U26660 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20840) );
  INV_X1 U26662 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20838) );
  INV_X1 U26664 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20835) );
  INV_X1 U26666 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20833) );
  INV_X1 U26668 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20832) );
  INV_X1 U26670 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20830) );
  INV_X1 U26672 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20827) );
  INV_X1 U26674 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20825) );
  INV_X1 U26676 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20816) );
  INV_X1 U26678 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20814) );
  INV_X1 U26680 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20811) );
  INV_X1 U26682 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20809) );
  INV_X1 U26684 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20776) );
  INV_X1 U26686 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20774) );
  INV_X1 U26688 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20771) );
  INV_X1 U26690 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20769) );
  INV_X1 U26692 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20712) );
  INV_X1 U26694 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20710) );
  INV_X1 U26696 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20707) );
  INV_X1 U26698 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20705) );
  INV_X1 U26700 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20688) );
  INV_X1 U26702 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20686) );
  INV_X1 U26704 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20683) );
  INV_X1 U26706 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20681) );
  INV_X1 U26708 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20616) );
  INV_X1 U26710 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20614) );
  INV_X1 U26712 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20611) );
  INV_X1 U26714 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20609) );
  INV_X1 U26716 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20592) );
  INV_X1 U26718 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20590) );
  INV_X1 U26720 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20587) );
  INV_X1 U26722 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20585) );
  INV_X1 U26724 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20536) );
  INV_X1 U26726 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20534) );
  INV_X1 U26728 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20531) );
  INV_X1 U26730 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20529) );
  INV_X1 U26732 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20528) );
  INV_X1 U26734 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20526) );
  INV_X1 U26736 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20523) );
  INV_X1 U26738 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20521) );
  INV_X1 U26740 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20392) );
  INV_X1 U26742 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20390) );
  INV_X1 U26744 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20387) );
  INV_X1 U26746 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20385) );
  INV_X1 U26748 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20384) );
  INV_X1 U26750 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20382) );
  INV_X1 U26752 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20379) );
  INV_X1 U26754 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20377) );
  INV_X1 U26756 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20280) );
  INV_X1 U26758 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20278) );
  INV_X1 U26760 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20275) );
  INV_X1 U26762 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20273) );
  INV_X1 U26764 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20264) );
  INV_X1 U26766 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20262) );
  INV_X1 U26768 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20259) );
  INV_X1 U26770 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20257) );
  INV_X1 U26772 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20216) );
  INV_X1 U26774 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20214) );
  INV_X1 U26776 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20211) );
  INV_X1 U26778 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20209) );
  INV_X1 U26780 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20184) );
  INV_X1 U26782 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20182) );
  INV_X1 U26784 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20179) );
  INV_X1 U26786 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20177) );
  INV_X1 U26788 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20160) );
  INV_X1 U26790 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20158) );
  INV_X1 U26792 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20155) );
  INV_X1 U26794 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20153) );
  INV_X1 U26796 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20120) );
  INV_X1 U26798 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20118) );
  INV_X1 U26800 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20115) );
  INV_X1 U26802 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20113) );
  INV_X1 U26804 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20103) );
  INV_X1 U26806 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20101) );
  INV_X1 U26808 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20100) );
  INV_X1 U26810 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20098) );
  INV_X1 U26812 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20096) );
  INV_X1 U26814 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20094) );
  INV_X1 U26816 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20091) );
  INV_X1 U26818 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20089) );
  INV_X1 U26820 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20088) );
  INV_X1 U26822 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20086) );
  INV_X1 U26824 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20083) );
  INV_X1 U26826 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20081) );
  INV_X1 U26828 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20064) );
  INV_X1 U26830 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20062) );
  INV_X1 U26832 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20059) );
  INV_X1 U26834 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20057) );
  INV_X1 U26836 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20056) );
  INV_X1 U26838 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20054) );
  INV_X1 U26840 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20051) );
  INV_X1 U26842 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20049) );
  INV_X1 U26844 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20048) );
  INV_X1 U26846 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20046) );
  INV_X1 U26848 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20043) );
  INV_X1 U26850 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20041) );
  INV_X1 U26852 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20032) );
  INV_X1 U26854 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20030) );
  INV_X1 U26856 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20027) );
  INV_X1 U26858 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20025) );
  INV_X1 U26860 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20016) );
  INV_X1 U26862 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20014) );
  INV_X1 U26864 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20011) );
  INV_X1 U26866 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20009) );
  INV_X1 U26868 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n20000) );
  INV_X1 U26870 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19998) );
  INV_X1 U26872 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19995) );
  INV_X1 U26874 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19993) );
  INV_X1 U26876 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19992) );
  INV_X1 U26878 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19990) );
  INV_X1 U26880 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19987) );
  INV_X1 U26882 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19985) );
  INV_X1 U26884 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19975) );
  INV_X1 U26886 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19973) );
  INV_X1 U26888 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19972) );
  INV_X1 U26890 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19970) );
  INV_X1 U26892 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19967) );
  INV_X1 U26894 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19965) );
  INV_X1 U26896 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19964) );
  INV_X1 U26898 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19962) );
  INV_X1 U26900 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19936) );
  INV_X1 U26902 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19934) );
  INV_X1 U26904 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19931) );
  INV_X1 U26906 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19929) );
  INV_X1 U26908 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19216) );
  INV_X1 U26910 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19214) );
  INV_X1 U26912 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19211) );
  INV_X1 U26914 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19209) );
  INV_X1 U26916 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19167) );
  INV_X1 U26918 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19165) );
  INV_X1 U26920 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19164) );
  INV_X1 U26922 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19162) );
  INV_X1 U26924 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19120) );
  INV_X1 U26926 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19118) );
  INV_X1 U26928 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19115) );
  INV_X1 U26930 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19113) );
  INV_X1 U26932 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19064) );
  INV_X1 U26934 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19062) );
  INV_X1 U26936 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19059) );
  INV_X1 U26938 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n19057) );
  INV_X1 U26940 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18992) );
  INV_X1 U26942 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18990) );
  INV_X1 U26944 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18987) );
  INV_X1 U26946 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18985) );
  INV_X1 U26948 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18928) );
  INV_X1 U26950 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18926) );
  INV_X1 U26952 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18923) );
  INV_X1 U26954 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18921) );
  INV_X1 U26956 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18880) );
  INV_X1 U26958 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18878) );
  INV_X1 U26960 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18875) );
  INV_X1 U26962 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18873) );
  INV_X1 U26964 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18856) );
  INV_X1 U26966 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18854) );
  INV_X1 U26968 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18851) );
  INV_X1 U26970 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18849) );
  INV_X1 U26972 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18792) );
  INV_X1 U26974 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18790) );
  INV_X1 U26976 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18787) );
  INV_X1 U26978 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18785) );
  INV_X1 U26980 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18784) );
  INV_X1 U26982 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18782) );
  INV_X1 U26984 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18779) );
  INV_X1 U26986 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18777) );
  INV_X1 U26988 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18768) );
  INV_X1 U26990 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18766) );
  INV_X1 U26992 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18763) );
  INV_X1 U26994 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18761) );
  INV_X1 U26996 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18728) );
  INV_X1 U26998 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18726) );
  INV_X1 U27000 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18723) );
  INV_X1 U27002 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18721) );
  INV_X1 U27004 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18664) );
  INV_X1 U27006 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18662) );
  INV_X1 U27008 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18659) );
  INV_X1 U27010 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18657) );
  INV_X1 U27012 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18640) );
  INV_X1 U27014 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18638) );
  INV_X1 U27016 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18635) );
  INV_X1 U27018 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18633) );
  INV_X1 U27020 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18568) );
  INV_X1 U27022 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18566) );
  INV_X1 U27024 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18563) );
  INV_X1 U27026 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18561) );
  INV_X1 U27028 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18544) );
  INV_X1 U27030 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18542) );
  INV_X1 U27032 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18539) );
  INV_X1 U27034 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18537) );
  INV_X1 U27036 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18488) );
  INV_X1 U27038 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18486) );
  INV_X1 U27040 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18483) );
  INV_X1 U27042 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18481) );
  INV_X1 U27044 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18480) );
  INV_X1 U27046 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18478) );
  INV_X1 U27048 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18475) );
  INV_X1 U27050 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18473) );
  INV_X1 U27052 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18344) );
  INV_X1 U27054 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18342) );
  INV_X1 U27056 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18339) );
  INV_X1 U27058 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18337) );
  INV_X1 U27060 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18336) );
  INV_X1 U27062 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18334) );
  INV_X1 U27064 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18331) );
  INV_X1 U27066 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18329) );
  INV_X1 U27068 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18232) );
  INV_X1 U27070 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18230) );
  INV_X1 U27072 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18227) );
  INV_X1 U27074 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18225) );
  INV_X1 U27076 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18216) );
  INV_X1 U27078 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18214) );
  INV_X1 U27080 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18211) );
  INV_X1 U27082 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18209) );
  INV_X1 U27084 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18168) );
  INV_X1 U27086 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18166) );
  INV_X1 U27088 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18163) );
  INV_X1 U27090 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18161) );
  INV_X1 U27092 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18136) );
  INV_X1 U27094 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18134) );
  INV_X1 U27096 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18131) );
  INV_X1 U27098 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18129) );
  INV_X1 U27100 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18112) );
  INV_X1 U27102 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18110) );
  INV_X1 U27104 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18107) );
  INV_X1 U27106 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18105) );
  INV_X1 U27108 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18072) );
  INV_X1 U27110 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18070) );
  INV_X1 U27112 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18067) );
  INV_X1 U27114 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18065) );
  INV_X1 U27116 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18055) );
  INV_X1 U27118 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18053) );
  INV_X1 U27120 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18052) );
  INV_X1 U27122 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18050) );
  INV_X1 U27124 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18048) );
  INV_X1 U27126 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18046) );
  INV_X1 U27128 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18043) );
  INV_X1 U27130 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18041) );
  INV_X1 U27132 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18040) );
  INV_X1 U27134 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18038) );
  INV_X1 U27136 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18035) );
  INV_X1 U27138 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18033) );
  INV_X1 U27140 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18016) );
  INV_X1 U27142 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18014) );
  INV_X1 U27144 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18011) );
  INV_X1 U27146 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18009) );
  INV_X1 U27148 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18008) );
  INV_X1 U27150 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18006) );
  INV_X1 U27152 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18003) );
  INV_X1 U27154 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18001) );
  INV_X1 U27156 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n18000) );
  INV_X1 U27158 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17998) );
  INV_X1 U27160 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17995) );
  INV_X1 U27162 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17993) );
  INV_X1 U27164 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17984) );
  INV_X1 U27166 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17982) );
  INV_X1 U27168 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17979) );
  INV_X1 U27170 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17977) );
  INV_X1 U27172 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17968) );
  INV_X1 U27174 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17966) );
  INV_X1 U27176 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17963) );
  INV_X1 U27178 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17961) );
  INV_X1 U27180 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17952) );
  INV_X1 U27182 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17950) );
  INV_X1 U27184 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17947) );
  INV_X1 U27186 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17945) );
  INV_X1 U27188 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17944) );
  INV_X1 U27190 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17942) );
  INV_X1 U27192 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17939) );
  INV_X1 U27194 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17937) );
  INV_X1 U27196 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17927) );
  INV_X1 U27198 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17925) );
  INV_X1 U27200 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17924) );
  INV_X1 U27202 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17922) );
  INV_X1 U27204 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17919) );
  INV_X1 U27206 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17917) );
  INV_X1 U27208 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17916) );
  INV_X1 U27210 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17914) );
  INV_X1 U27212 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17888) );
  INV_X1 U27214 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17886) );
  INV_X1 U27216 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17883) );
  INV_X1 U27218 ( .A(1'b1), .ZN(p_wishbone_bd_ram_n17881) );
  INV_X1 U27220 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n185) );
  INV_X1 U27222 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n184) );
  INV_X1 U27224 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n181) );
  INV_X1 U27226 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n182) );
  INV_X1 U27228 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n183) );
  INV_X1 U27230 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n180) );
  INV_X1 U27232 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n179) );
  INV_X1 U27234 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n177) );
  INV_X1 U27236 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n178) );
  INV_X1 U27238 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n161) );
  INV_X1 U27240 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n176) );
  INV_X1 U27242 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n162) );
  INV_X1 U27244 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n163) );
  INV_X1 U27246 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n164) );
  INV_X1 U27248 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n165) );
  INV_X1 U27250 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n166) );
  INV_X1 U27252 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n167) );
  INV_X1 U27254 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n168) );
  INV_X1 U27256 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n169) );
  INV_X1 U27258 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n170) );
  INV_X1 U27260 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n171) );
  INV_X1 U27262 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n172) );
  INV_X1 U27264 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n173) );
  INV_X1 U27266 ( .A(1'b1), .ZN(p_rxethmac1_rxcounters1_n174) );
  INV_X1 U27268 ( .A(1'b0), .ZN(p_rxethmac1_rxcounters1_n175) );
  INV_X1 U27270 ( .A(1'b1), .ZN(p_rxethmac1_rxstatem1_n40) );
  INV_X1 U27272 ( .A(1'b0), .ZN(p_rxethmac1_rxstatem1_n38) );
  INV_X1 U27274 ( .A(1'b0), .ZN(p_txethmac1_random1_n108) );
  INV_X1 U27276 ( .A(1'b1), .ZN(p_txethmac1_random1_x_0) );
  INV_X1 U27278 ( .A(1'b1), .ZN(p_txethmac1_random1_x_1) );
  INV_X1 U27280 ( .A(1'b1), .ZN(p_txethmac1_random1_x_2) );
  INV_X1 U27282 ( .A(1'b1), .ZN(p_txethmac1_random1_x_3) );
  INV_X1 U27284 ( .A(1'b1), .ZN(p_txethmac1_random1_x_4) );
  INV_X1 U27286 ( .A(1'b1), .ZN(p_txethmac1_random1_x_5) );
  INV_X1 U27288 ( .A(1'b1), .ZN(p_txethmac1_random1_x_6) );
  INV_X1 U27290 ( .A(1'b1), .ZN(p_txethmac1_random1_x_7) );
  INV_X1 U27292 ( .A(1'b1), .ZN(p_txethmac1_random1_x_8) );
  INV_X1 U27294 ( .A(1'b0), .ZN(p_txethmac1_random1_n107) );
  INV_X1 U27296 ( .A(1'b1), .ZN(p_txethmac1_random1_n106) );
  INV_X1 U27298 ( .A(1'b1), .ZN(p_txethmac1_random1_n105) );
  INV_X1 U27300 ( .A(1'b0), .ZN(p_txethmac1_random1_n104) );
  INV_X1 U27302 ( .A(1'b0), .ZN(p_txethmac1_random1_n103) );
  INV_X1 U27304 ( .A(1'b0), .ZN(p_txethmac1_random1_n102) );
  INV_X1 U27306 ( .A(1'b0), .ZN(p_txethmac1_random1_n101) );
  INV_X1 U27308 ( .A(1'b1), .ZN(p_txethmac1_random1_n100) );
  INV_X1 U27310 ( .A(1'b0), .ZN(p_txethmac1_random1_n99) );
  INV_X1 U27312 ( .A(1'b1), .ZN(p_txethmac1_random1_n98) );
  INV_X1 U27314 ( .A(1'b0), .ZN(p_txethmac1_txcrc_N27) );
  INV_X1 U27316 ( .A(1'b0), .ZN(p_txethmac1_txcrc_N12) );
  INV_X1 U27318 ( .A(1'b1), .ZN(p_txethmac1_txcrc_N4) );
  INV_X1 U27320 ( .A(1'b0), .ZN(p_txethmac1_txcrc_N9) );
  INV_X1 U27322 ( .A(1'b0), .ZN(p_txethmac1_txstatem1_n92) );
  INV_X1 U27324 ( .A(1'b1), .ZN(p_txethmac1_StateJam) );
  INV_X1 U27326 ( .A(1'b0), .ZN(p_txethmac1_txstatem1_n90) );
  INV_X1 U27328 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n206) );
  INV_X1 U27330 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n205) );
  INV_X1 U27332 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n203) );
  INV_X1 U27334 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n204) );
  INV_X1 U27336 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n202) );
  INV_X1 U27338 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n201) );
  INV_X1 U27340 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n200) );
  INV_X1 U27342 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n199) );
  INV_X1 U27344 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n198) );
  INV_X1 U27346 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n197) );
  INV_X1 U27348 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n196) );
  INV_X1 U27350 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n195) );
  INV_X1 U27352 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n194) );
  INV_X1 U27354 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n192) );
  INV_X1 U27356 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n191) );
  INV_X1 U27358 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n190) );
  INV_X1 U27360 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n189) );
  INV_X1 U27362 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n175) );
  INV_X1 U27364 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n176) );
  INV_X1 U27366 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n177) );
  INV_X1 U27368 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n178) );
  INV_X1 U27370 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n179) );
  INV_X1 U27372 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n180) );
  INV_X1 U27374 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n181) );
  INV_X1 U27376 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n182) );
  INV_X1 U27378 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n183) );
  INV_X1 U27380 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n184) );
  INV_X1 U27382 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n185) );
  INV_X1 U27384 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n186) );
  INV_X1 U27386 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n187) );
  INV_X1 U27388 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n188) );
  INV_X1 U27390 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n174) );
  INV_X1 U27392 ( .A(1'b0), .ZN(p_txethmac1_txcounters1_n173) );
  INV_X1 U27394 ( .A(1'b1), .ZN(p_txethmac1_txcounters1_n172) );
  INV_X1 U27396 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n284) );
  INV_X1 U27398 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n281) );
  INV_X1 U27400 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n280) );
  INV_X1 U27402 ( .A(1'b1), .ZN(p_maccontrol1_TxCtrlStartFrm) );
  INV_X1 U27404 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n271) );
  INV_X1 U27406 ( .A(1'b1), .ZN(p_maccontrol1_transmitcontrol1_n278) );
  INV_X1 U27408 ( .A(1'b1), .ZN(p_maccontrol1_transmitcontrol1_n277) );
  INV_X1 U27410 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n283) );
  INV_X1 U27412 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n272) );
  INV_X1 U27414 ( .A(1'b0), .ZN(p_maccontrol1_transmitcontrol1_n275) );
  INV_X1 U27416 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n570) );
  INV_X1 U27418 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n568) );
  INV_X1 U27420 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n567) );
  INV_X1 U27422 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n566) );
  INV_X1 U27424 ( .A(1'b1), .ZN(p_maccontrol1_receivecontrol1_n562) );
  INV_X1 U27426 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n563) );
  INV_X1 U27428 ( .A(1'b1), .ZN(p_maccontrol1_receivecontrol1_n564) );
  INV_X1 U27430 ( .A(1'b1), .ZN(p_maccontrol1_receivecontrol1_n560) );
  INV_X1 U27432 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n525) );
  INV_X1 U27434 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n524) );
  INV_X1 U27436 ( .A(1'b1), .ZN(p_maccontrol1_receivecontrol1_n504) );
  INV_X1 U27438 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n505) );
  INV_X1 U27440 ( .A(1'b1), .ZN(p_maccontrol1_receivecontrol1_n506) );
  INV_X1 U27442 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n507) );
  INV_X1 U27444 ( .A(1'b0), .ZN(p_maccontrol1_receivecontrol1_n503) );
  INV_X1 U27446 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n52) );
  INV_X1 U27448 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n51) );
  INV_X1 U27450 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n50) );
  INV_X1 U27452 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n49) );
  INV_X1 U27454 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n48) );
  INV_X1 U27456 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n47) );
  INV_X1 U27458 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n46) );
  INV_X1 U27460 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n45) );
  INV_X1 U27462 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n44) );
  INV_X1 U27464 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n43) );
  INV_X1 U27466 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n42) );
  INV_X1 U27468 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n41) );
  INV_X1 U27470 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n40) );
  INV_X1 U27472 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n39) );
  INV_X1 U27474 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n38) );
  INV_X1 U27476 ( .A(1'b0), .ZN(p_ethreg1_MIIRX_DATA_n37) );
  INV_X1 U27478 ( .A(1'b0), .ZN(p_ethreg1_MIIADDRESS_0_n19) );
  INV_X1 U27480 ( .A(1'b0), .ZN(p_ethreg1_MIIADDRESS_0_n18) );
  INV_X1 U27482 ( .A(1'b0), .ZN(p_ethreg1_MIIADDRESS_0_n17) );
  INV_X1 U27484 ( .A(1'b0), .ZN(p_ethreg1_MIIADDRESS_0_n16) );
  INV_X1 U27486 ( .A(1'b0), .ZN(p_ethreg1_MIIADDRESS_0_n15) );
  INV_X1 U27488 ( .A(1'b0), .ZN(n33932) );
  INV_X1 U27490 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n31) );
  INV_X1 U27492 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n30) );
  INV_X1 U27494 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n29) );
  INV_X1 U27496 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n28) );
  INV_X1 U27498 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n27) );
  INV_X1 U27500 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n26) );
  INV_X1 U27502 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n25) );
  INV_X1 U27504 ( .A(1'b0), .ZN(p_ethreg1_MIIMODER_0_n24) );
  INV_X1 U27506 ( .A(1'b0), .ZN(p_ethreg1_CTRLMODER_0_n12) );
  INV_X1 U27508 ( .A(1'b0), .ZN(p_ethreg1_CTRLMODER_0_n11) );
  INV_X1 U27510 ( .A(1'b0), .ZN(p_ethreg1_CTRLMODER_0_n10) );
  INV_X1 U27512 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_2_n18) );
  INV_X1 U27514 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_2_n17) );
  INV_X1 U27516 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_2_n16) );
  INV_X1 U27518 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_2_n15) );
  INV_X1 U27520 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n26) );
  INV_X1 U27522 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n25) );
  INV_X1 U27524 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n24) );
  INV_X1 U27526 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n23) );
  INV_X1 U27528 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n22) );
  INV_X1 U27530 ( .A(1'b0), .ZN(p_ethreg1_COLLCONF_0_n21) );
  INV_X1 U27532 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n29) );
  INV_X1 U27534 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n17) );
  INV_X1 U27536 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n27) );
  INV_X1 U27538 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n26) );
  INV_X1 U27540 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n25) );
  INV_X1 U27542 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n24) );
  INV_X1 U27544 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n23) );
  INV_X1 U27546 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_2_n22) );
  INV_X1 U27548 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n30) );
  INV_X1 U27550 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n29) );
  INV_X1 U27552 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n28) );
  INV_X1 U27554 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n27) );
  INV_X1 U27556 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n26) );
  INV_X1 U27558 ( .A(1'b0), .ZN(n33923) );
  INV_X1 U27560 ( .A(1'b0), .ZN(n33924) );
  INV_X1 U27562 ( .A(1'b0), .ZN(p_ethreg1_PACKETLEN_1_n23) );
  INV_X1 U27564 ( .A(1'b0), .ZN(p_ethreg1_IPGR1_0_n27) );
  INV_X1 U27566 ( .A(1'b0), .ZN(p_ethreg1_IPGR1_0_n26) );
  INV_X1 U27568 ( .A(1'b0), .ZN(p_ethreg1_IPGR1_0_n25) );
  INV_X1 U27570 ( .A(1'b0), .ZN(n33928) );
  INV_X1 U27572 ( .A(1'b0), .ZN(n33929) );
  INV_X1 U27574 ( .A(1'b0), .ZN(p_ethreg1_IPGR1_0_n22) );
  INV_X1 U27576 ( .A(1'b0), .ZN(p_ethreg1_IPGR1_0_n21) );
  INV_X1 U27578 ( .A(1'b0), .ZN(p_ethreg1_IPGT_0_n27) );
  INV_X1 U27580 ( .A(1'b0), .ZN(p_ethreg1_IPGT_0_n26) );
  INV_X1 U27582 ( .A(1'b0), .ZN(n33927) );
  INV_X1 U27584 ( .A(1'b0), .ZN(p_ethreg1_IPGT_0_n24) );
  INV_X1 U27586 ( .A(1'b0), .ZN(p_ethreg1_IPGT_0_n23) );
  INV_X1 U27588 ( .A(1'b0), .ZN(n33931) );
  INV_X1 U27590 ( .A(1'b0), .ZN(p_ethreg1_IPGT_0_n21) );
  INV_X1 U27592 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n25) );
  INV_X1 U27594 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n24) );
  INV_X1 U27596 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n23) );
  INV_X1 U27598 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n22) );
  INV_X1 U27600 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n21) );
  INV_X1 U27602 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n20) );
  INV_X1 U27604 ( .A(1'b0), .ZN(p_ethreg1_INT_MASK_0_n19) );
  INV_X1 U27606 ( .A(1'b0), .ZN(n33921) );
  INV_X1 U27608 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n29) );
  INV_X1 U27610 ( .A(1'b0), .ZN(n33922) );
  INV_X1 U27612 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n27) );
  INV_X1 U27614 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n26) );
  INV_X1 U27616 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n25) );
  INV_X1 U27618 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n24) );
  INV_X1 U27620 ( .A(1'b0), .ZN(p_ethreg1_MODER_1_n23) );
  INV_X1 U27622 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n28) );
  INV_X1 U27624 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n27) );
  INV_X1 U27626 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n26) );
  INV_X1 U27628 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n25) );
  INV_X1 U27630 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n24) );
  INV_X1 U27632 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n23) );
  INV_X1 U27634 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n22) );
  INV_X1 U27636 ( .A(1'b0), .ZN(p_ethreg1_MODER_0_n21) );
  INV_X1 U27638 ( .A(1'b1), .ZN(p_miim1_outctrl_n36) );
  INV_X1 U27640 ( .A(1'b1), .ZN(p_miim1_outctrl_n35) );
  INV_X1 U27642 ( .A(1'b1), .ZN(p_miim1_outctrl_n33) );
  INV_X1 U27644 ( .A(1'b0), .ZN(p_miim1_shftrg_n161) );
  INV_X1 U27646 ( .A(1'b0), .ZN(p_miim1_shftrg_n160) );
  INV_X1 U27648 ( .A(1'b0), .ZN(p_miim1_shftrg_n159) );
  INV_X1 U27650 ( .A(1'b0), .ZN(p_miim1_shftrg_n158) );
  INV_X1 U27652 ( .A(1'b0), .ZN(p_miim1_shftrg_n157) );
  INV_X1 U27654 ( .A(1'b0), .ZN(p_miim1_shftrg_n156) );
  INV_X1 U27656 ( .A(1'b0), .ZN(p_miim1_shftrg_n155) );
  INV_X1 U27658 ( .A(1'b0), .ZN(p_miim1_shftrg_n154) );
  INV_X1 U27660 ( .A(1'b0), .ZN(p_miim1_shftrg_n153) );
  INV_X1 U27662 ( .A(1'b0), .ZN(p_miim1_shftrg_n152) );
  INV_X1 U27664 ( .A(1'b0), .ZN(p_miim1_shftrg_n151) );
  INV_X1 U27666 ( .A(1'b0), .ZN(p_miim1_shftrg_n150) );
  INV_X1 U27668 ( .A(1'b0), .ZN(p_miim1_shftrg_n149) );
  INV_X1 U27670 ( .A(1'b0), .ZN(p_miim1_shftrg_n148) );
  INV_X1 U27672 ( .A(1'b0), .ZN(p_miim1_shftrg_n147) );
  INV_X1 U27674 ( .A(1'b0), .ZN(p_miim1_shftrg_n146) );
  INV_X1 U27676 ( .A(1'b0), .ZN(p_miim1_clkgen_N15) );
  INV_X1 U27678 ( .A(1'b0), .ZN(p_miim1_clkgen_N16) );
  INV_X1 U27680 ( .A(1'b0), .ZN(p_miim1_clkgen_N17) );
  INV_X1 U27682 ( .A(1'b0), .ZN(p_miim1_clkgen_N18) );
  INV_X1 U27684 ( .A(1'b0), .ZN(p_miim1_clkgen_N19) );
  INV_X1 U27686 ( .A(1'b0), .ZN(p_miim1_clkgen_N20) );
  INV_X1 U27688 ( .A(1'b0), .ZN(p_miim1_clkgen_N21) );
  INV_X1 U27690 ( .A(1'b1), .ZN(p_miim1_clkgen_n35) );
  INV_X1 U27692 ( .A(1'b0), .ZN(p_macstatus1_n97) );
  INV_X1 U27694 ( .A(1'b0), .ZN(p_macstatus1_N7) );
  INV_X1 U27696 ( .A(1'b1), .ZN(p_macstatus1_TakeSample) );
  INV_X1 U27698 ( .A(1'b1), .ZN(LoadRxStatus) );
  INV_X1 U27700 ( .A(1'b0), .ZN(p_macstatus1_n95) );
  INV_X1 U27702 ( .A(1'b0), .ZN(p_macstatus1_n93) );
  INV_X1 U27704 ( .A(1'b0), .ZN(p_macstatus1_n91) );
  INV_X1 U27706 ( .A(1'b0), .ZN(p_macstatus1_n87) );
  INV_X1 U27708 ( .A(1'b0), .ZN(p_macstatus1_n86) );
  INV_X1 U27710 ( .A(1'b0), .ZN(p_macstatus1_n85) );
  INV_X1 U27712 ( .A(1'b0), .ZN(p_macstatus1_n84) );
  INV_X1 U27714 ( .A(1'b0), .ZN(p_macstatus1_n90) );
  INV_X1 U27716 ( .A(1'b0), .ZN(p_wishbone_n2474) );
  INV_X1 U27718 ( .A(1'b1), .ZN(p_wishbone_TxRetry_wb) );
  INV_X1 U27720 ( .A(1'b1), .ZN(p_wishbone_TxDone_wb) );
  INV_X1 U27722 ( .A(1'b1), .ZN(p_wishbone_TxAbort_wb) );
  INV_X1 U27724 ( .A(1'b1), .ZN(p_wishbone_LatchedRxStartFrm) );
  INV_X1 U27726 ( .A(1'b1), .ZN(p_wishbone_SyncRxStartFrm_q) );
  INV_X1 U27728 ( .A(1'b1), .ZN(p_wishbone_RxAbortLatched) );
  INV_X1 U27730 ( .A(1'b1), .ZN(p_wishbone_RxAbortSync3) );
  INV_X1 U27732 ( .A(1'b1), .ZN(p_wishbone_RxAbortSync2) );
  INV_X1 U27734 ( .A(1'b0), .ZN(p_wishbone_n2133) );
  INV_X1 U27736 ( .A(1'b0), .ZN(p_wishbone_n2132) );
  INV_X1 U27738 ( .A(1'b0), .ZN(p_wishbone_n2131) );
  INV_X1 U27740 ( .A(1'b0), .ZN(p_wishbone_n2130) );
  INV_X1 U27742 ( .A(1'b0), .ZN(p_wishbone_n2129) );
  INV_X1 U27744 ( .A(1'b0), .ZN(p_wishbone_n2128) );
  INV_X1 U27746 ( .A(1'b0), .ZN(p_wishbone_n2127) );
  INV_X1 U27748 ( .A(1'b0), .ZN(p_wishbone_n2126) );
  INV_X1 U27750 ( .A(1'b0), .ZN(p_wishbone_n2125) );
  INV_X1 U27752 ( .A(1'b0), .ZN(p_wishbone_n2124) );
  INV_X1 U27754 ( .A(1'b0), .ZN(p_wishbone_n2123) );
  INV_X1 U27756 ( .A(1'b0), .ZN(p_wishbone_n2122) );
  INV_X1 U27758 ( .A(1'b0), .ZN(p_wishbone_n2121) );
  INV_X1 U27760 ( .A(1'b0), .ZN(p_wishbone_n2120) );
  INV_X1 U27762 ( .A(1'b0), .ZN(p_wishbone_n2119) );
  INV_X1 U27764 ( .A(1'b0), .ZN(p_wishbone_n2118) );
  INV_X1 U27766 ( .A(1'b0), .ZN(p_wishbone_n2117) );
  INV_X1 U27768 ( .A(1'b0), .ZN(p_wishbone_n2115) );
  INV_X1 U27770 ( .A(1'b0), .ZN(p_wishbone_n2112) );
  INV_X1 U27772 ( .A(1'b0), .ZN(p_wishbone_n2111) );
  INV_X1 U27774 ( .A(1'b1), .ZN(p_wishbone_LatchValidBytes) );
  INV_X1 U27776 ( .A(1'b1), .ZN(p_wishbone_n2300) );
  INV_X1 U27778 ( .A(1'b1), .ZN(p_wishbone_n2298) );
  INV_X1 U27780 ( .A(1'b1), .ZN(p_wishbone_n2296) );
  INV_X1 U27782 ( .A(1'b1), .ZN(p_wishbone_ReadTxDataFromFifo_tck) );
  INV_X1 U27784 ( .A(1'b1), .ZN(p_wishbone_ReadTxDataFromFifo_syncb2) );
  INV_X1 U27786 ( .A(1'b1), .ZN(p_wishbone_ReadTxDataFromFifo_sync2) );
  INV_X1 U27788 ( .A(1'b0), .ZN(p_wishbone_n2465) );
  INV_X1 U27790 ( .A(1'b1), .ZN(p_wishbone_n2464) );
  INV_X1 U27792 ( .A(1'b1), .ZN(p_wishbone_n2466) );
  INV_X1 U27794 ( .A(1'b1), .ZN(p_wishbone_n2346) );
  INV_X1 U27796 ( .A(1'b0), .ZN(p_wishbone_n2345) );
  INV_X1 U27798 ( .A(1'b1), .ZN(p_wishbone_n2344) );
  INV_X1 U27800 ( .A(1'b0), .ZN(p_wishbone_n2343) );
  INV_X1 U27802 ( .A(1'b1), .ZN(p_wishbone_n2463) );
  INV_X1 U27804 ( .A(1'b0), .ZN(n33934) );
  INV_X1 U27806 ( .A(1'b1), .ZN(p_wishbone_N867) );
  INV_X1 U27808 ( .A(1'b0), .ZN(p_wishbone_n2461) );
  INV_X1 U27810 ( .A(1'b1), .ZN(p_wishbone_n2317) );
  INV_X1 U27812 ( .A(1'b1), .ZN(p_wishbone_n2318) );
  INV_X1 U27814 ( .A(1'b0), .ZN(p_wishbone_n2457) );
  INV_X1 U27816 ( .A(1'b1), .ZN(p_wishbone_TxEn) );
  INV_X1 U27818 ( .A(1'b0), .ZN(p_wishbone_n2319) );
  INV_X1 U27820 ( .A(1'b0), .ZN(p_wishbone_n2108) );
  INV_X1 U27822 ( .A(1'b0), .ZN(p_wishbone_n2107) );
  INV_X1 U27824 ( .A(1'b0), .ZN(p_wishbone_n2106) );
  INV_X1 U27826 ( .A(1'b0), .ZN(p_wishbone_n2105) );
  INV_X1 U27828 ( .A(1'b1), .ZN(p_wishbone_n2299) );
  INV_X1 U27830 ( .A(1'b1), .ZN(p_wishbone_n2320) );
  INV_X1 U27832 ( .A(1'b0), .ZN(p_wishbone_n2104) );
  INV_X1 U27834 ( .A(1'b0), .ZN(p_wishbone_n2103) );
  INV_X1 U27836 ( .A(1'b0), .ZN(p_wishbone_n2102) );
  INV_X1 U27838 ( .A(1'b0), .ZN(p_wishbone_n2101) );
  INV_X1 U27840 ( .A(1'b0), .ZN(p_wishbone_n2100) );
  INV_X1 U27842 ( .A(1'b0), .ZN(p_wishbone_n2099) );
  INV_X1 U27844 ( .A(1'b0), .ZN(p_wishbone_n2098) );
  INV_X1 U27846 ( .A(1'b0), .ZN(p_wishbone_n2097) );
  INV_X1 U27848 ( .A(1'b0), .ZN(p_wishbone_n2096) );
  INV_X1 U27850 ( .A(1'b0), .ZN(p_wishbone_n2095) );
  INV_X1 U27852 ( .A(1'b0), .ZN(p_wishbone_n2094) );
  INV_X1 U27854 ( .A(1'b0), .ZN(p_wishbone_n2093) );
  INV_X1 U27856 ( .A(1'b0), .ZN(p_wishbone_n2092) );
  INV_X1 U27858 ( .A(1'b0), .ZN(p_wishbone_n2091) );
  INV_X1 U27860 ( .A(1'b0), .ZN(p_wishbone_n2090) );
  INV_X1 U27862 ( .A(1'b0), .ZN(p_wishbone_n2089) );
  INV_X1 U27864 ( .A(1'b1), .ZN(p_wishbone_n2330) );
  INV_X1 U27866 ( .A(1'b1), .ZN(p_wishbone_WbEn) );
  INV_X1 U27868 ( .A(1'b0), .ZN(p_wishbone_n2428) );
  INV_X1 U27870 ( .A(1'b1), .ZN(p_wishbone_RxEn) );
  INV_X1 U27872 ( .A(1'b0), .ZN(p_wishbone_n2326) );
  INV_X1 U27874 ( .A(1'b0), .ZN(p_wishbone_n2417) );
  INV_X1 U27876 ( .A(1'b0), .ZN(p_wishbone_n2415) );
  INV_X1 U27878 ( .A(1'b0), .ZN(p_wishbone_n2416) );
  INV_X1 U27880 ( .A(1'b0), .ZN(p_wishbone_n2391) );
  INV_X1 U27882 ( .A(1'b0), .ZN(p_wishbone_n2392) );
  INV_X1 U27884 ( .A(1'b0), .ZN(p_wishbone_n2393) );
  INV_X1 U27886 ( .A(1'b0), .ZN(p_wishbone_n2394) );
  INV_X1 U27888 ( .A(1'b0), .ZN(p_wishbone_n2395) );
  INV_X1 U27890 ( .A(1'b0), .ZN(p_wishbone_n2396) );
  INV_X1 U27892 ( .A(1'b0), .ZN(p_wishbone_n2397) );
  INV_X1 U27894 ( .A(1'b0), .ZN(p_wishbone_n2398) );
  INV_X1 U27896 ( .A(1'b0), .ZN(p_wishbone_n2425) );
  INV_X1 U27898 ( .A(1'b0), .ZN(p_wishbone_n2412) );
  INV_X1 U27900 ( .A(1'b1), .ZN(p_wishbone_ShiftEnded_rck) );
  INV_X1 U27902 ( .A(1'b1), .ZN(p_wishbone_ShiftEndedSync1) );
  INV_X1 U27904 ( .A(1'b1), .ZN(p_wishbone_ShiftEndedSync2) );
  INV_X1 U27906 ( .A(1'b1), .ZN(p_wishbone_ShiftEndedSync_c1) );
  INV_X1 U27908 ( .A(1'b0), .ZN(p_wishbone_n2413) );
  INV_X1 U27910 ( .A(1'b1), .ZN(p_wishbone_WriteRxDataToFifo) );
  INV_X1 U27912 ( .A(1'b1), .ZN(p_wishbone_WriteRxDataToFifoSync2) );
  INV_X1 U27914 ( .A(1'b0), .ZN(p_wishbone_n2383) );
  INV_X1 U27916 ( .A(1'b0), .ZN(p_wishbone_n2384) );
  INV_X1 U27918 ( .A(1'b0), .ZN(p_wishbone_n2385) );
  INV_X1 U27920 ( .A(1'b0), .ZN(p_wishbone_n2386) );
  INV_X1 U27922 ( .A(1'b0), .ZN(p_wishbone_n2387) );
  INV_X1 U27924 ( .A(1'b0), .ZN(p_wishbone_n2388) );
  INV_X1 U27926 ( .A(1'b0), .ZN(p_wishbone_n2389) );
  INV_X1 U27928 ( .A(1'b0), .ZN(p_wishbone_n2390) );
  INV_X1 U27930 ( .A(1'b0), .ZN(p_wishbone_n2352) );
  INV_X1 U27932 ( .A(1'b0), .ZN(p_wishbone_n2351) );
  INV_X1 U27934 ( .A(1'b0), .ZN(p_wishbone_n2354) );
  INV_X1 U27936 ( .A(1'b0), .ZN(p_wishbone_n2353) );
  INV_X1 U27938 ( .A(1'b0), .ZN(p_wishbone_n2356) );
  INV_X1 U27940 ( .A(1'b0), .ZN(p_wishbone_n2355) );
  INV_X1 U27942 ( .A(1'b0), .ZN(p_wishbone_n2358) );
  INV_X1 U27944 ( .A(1'b0), .ZN(p_wishbone_n2357) );
  INV_X1 U27946 ( .A(1'b0), .ZN(p_wishbone_n2360) );
  INV_X1 U27948 ( .A(1'b0), .ZN(p_wishbone_n2359) );
  INV_X1 U27950 ( .A(1'b0), .ZN(p_wishbone_n2362) );
  INV_X1 U27952 ( .A(1'b0), .ZN(p_wishbone_n2361) );
  INV_X1 U27954 ( .A(1'b0), .ZN(p_wishbone_n2364) );
  INV_X1 U27956 ( .A(1'b0), .ZN(p_wishbone_n2363) );
  INV_X1 U27958 ( .A(1'b0), .ZN(p_wishbone_n2366) );
  INV_X1 U27960 ( .A(1'b0), .ZN(p_wishbone_n2365) );
  INV_X1 U27962 ( .A(1'b0), .ZN(p_wishbone_n2399) );
  INV_X1 U27964 ( .A(1'b0), .ZN(p_wishbone_n2400) );
  INV_X1 U27966 ( .A(1'b0), .ZN(p_wishbone_n2401) );
  INV_X1 U27968 ( .A(1'b0), .ZN(p_wishbone_n2402) );
  INV_X1 U27970 ( .A(1'b0), .ZN(p_wishbone_n2403) );
  INV_X1 U27972 ( .A(1'b0), .ZN(p_wishbone_n2404) );
  INV_X1 U27974 ( .A(1'b0), .ZN(p_wishbone_n2405) );
  INV_X1 U27976 ( .A(1'b0), .ZN(p_wishbone_n2406) );
  INV_X1 U27978 ( .A(1'b0), .ZN(p_wishbone_n2325) );
  INV_X1 U27980 ( .A(1'b0), .ZN(p_wishbone_n2088) );
  INV_X1 U27982 ( .A(1'b0), .ZN(p_wishbone_n2087) );
  INV_X1 U27984 ( .A(1'b1), .ZN(p_wishbone_n2331) );
  INV_X1 U27986 ( .A(1'b0), .ZN(p_wishbone_n2247) );
  INV_X1 U27988 ( .A(1'b1), .ZN(p_wishbone_n2246) );
  INV_X1 U27990 ( .A(1'b0), .ZN(p_wishbone_n2245) );
  INV_X1 U27992 ( .A(1'b1), .ZN(p_wishbone_n2244) );
  INV_X1 U27994 ( .A(1'b0), .ZN(p_wishbone_n2243) );
  INV_X1 U27996 ( .A(1'b1), .ZN(p_wishbone_n2242) );
  INV_X1 U27998 ( .A(1'b0), .ZN(p_wishbone_n2241) );
  INV_X1 U28000 ( .A(1'b1), .ZN(p_wishbone_BlockingTxStatusWrite) );
  INV_X1 U28002 ( .A(1'b1), .ZN(p_wishbone_BlockingTxStatusWrite_sync2) );
  INV_X1 U28004 ( .A(1'b0), .ZN(n33933) );
  INV_X1 U28006 ( .A(1'b0), .ZN(p_wishbone_n2249) );
  INV_X1 U28008 ( .A(1'b0), .ZN(p_wishbone_n2294) );
  INV_X1 U28010 ( .A(1'b1), .ZN(p_wishbone_TxStartFrm_wb) );
  INV_X1 U28012 ( .A(1'b1), .ZN(p_wishbone_TxStartFrm_sync2) );
  INV_X1 U28014 ( .A(1'b1), .ZN(p_wishbone_n2291) );
  INV_X1 U28016 ( .A(1'b0), .ZN(p_wishbone_n2289) );
  INV_X1 U28018 ( .A(1'b0), .ZN(p_wishbone_n2288) );
  INV_X1 U28020 ( .A(1'b0), .ZN(p_wishbone_n2287) );
  INV_X1 U28022 ( .A(1'b0), .ZN(p_wishbone_n2286) );
  INV_X1 U28024 ( .A(1'b0), .ZN(p_wishbone_n2285) );
  INV_X1 U28026 ( .A(1'b0), .ZN(p_wishbone_n2284) );
  INV_X1 U28028 ( .A(1'b0), .ZN(p_wishbone_n2283) );
  INV_X1 U28030 ( .A(1'b0), .ZN(p_wishbone_n2282) );
  INV_X1 U28032 ( .A(1'b0), .ZN(p_wishbone_n2281) );
  INV_X1 U28034 ( .A(1'b0), .ZN(p_wishbone_n2280) );
  INV_X1 U28036 ( .A(1'b0), .ZN(p_wishbone_n2279) );
  INV_X1 U28038 ( .A(1'b0), .ZN(p_wishbone_n2278) );
  INV_X1 U28040 ( .A(1'b0), .ZN(p_wishbone_n2277) );
  INV_X1 U28042 ( .A(1'b0), .ZN(p_wishbone_n2276) );
  INV_X1 U28044 ( .A(1'b0), .ZN(p_wishbone_n2275) );
  INV_X1 U28046 ( .A(1'b0), .ZN(p_wishbone_n2274) );
  INV_X1 U28048 ( .A(1'b0), .ZN(p_wishbone_n2273) );
  INV_X1 U28050 ( .A(1'b0), .ZN(p_wishbone_n2272) );
  INV_X1 U28052 ( .A(1'b0), .ZN(p_wishbone_n2271) );
  INV_X1 U28054 ( .A(1'b0), .ZN(p_wishbone_n2270) );
  INV_X1 U28056 ( .A(1'b0), .ZN(p_wishbone_n2269) );
  INV_X1 U28058 ( .A(1'b0), .ZN(p_wishbone_n2268) );
  INV_X1 U28060 ( .A(1'b0), .ZN(p_wishbone_n2267) );
  INV_X1 U28062 ( .A(1'b0), .ZN(p_wishbone_n2266) );
  INV_X1 U28064 ( .A(1'b0), .ZN(p_wishbone_n2265) );
  INV_X1 U28066 ( .A(1'b0), .ZN(p_wishbone_n2264) );
  INV_X1 U28068 ( .A(1'b0), .ZN(p_wishbone_n2263) );
  INV_X1 U28070 ( .A(1'b0), .ZN(p_wishbone_n2262) );
  INV_X1 U28072 ( .A(1'b0), .ZN(p_wishbone_n2261) );
  INV_X1 U28074 ( .A(1'b0), .ZN(p_wishbone_n2260) );
  INV_X1 U28076 ( .A(1'b0), .ZN(p_wishbone_n2259) );
  INV_X1 U28078 ( .A(1'b0), .ZN(p_wishbone_n2258) );
  INV_X1 U28080 ( .A(1'b1), .ZN(p_wishbone_n2340) );
  INV_X1 U28082 ( .A(1'b1), .ZN(p_wishbone_n2341) );
  INV_X1 U28084 ( .A(1'b1), .ZN(p_wishbone_n2342) );
  INV_X1 U28086 ( .A(1'b1), .ZN(p_wishbone_n2339) );
  INV_X1 U28088 ( .A(1'b1), .ZN(p_wishbone_n2168) );
  INV_X1 U28090 ( .A(1'b1), .ZN(p_wishbone_n2141) );
  INV_X1 U28092 ( .A(1'b1), .ZN(p_wishbone_RxStatusWriteLatched) );
  INV_X1 U28094 ( .A(1'b1), .ZN(RxStatusWriteLatched_sync2) );
  INV_X1 U28096 ( .A(1'b0), .ZN(p_wishbone_n2138) );
  INV_X1 U28098 ( .A(1'b1), .ZN(p_wishbone_Busy_IRQ_rck) );
  INV_X1 U28100 ( .A(1'b1), .ZN(p_wishbone_Busy_IRQ_sync2) );
  INV_X1 U28102 ( .A(1'b0), .ZN(p_rxethmac1_N3) );
  INV_X1 U28104 ( .A(1'b1), .ZN(MRxD_Lb_3) );
  INV_X1 U28106 ( .A(1'b1), .ZN(MRxD_Lb_2) );
  INV_X1 U28108 ( .A(1'b1), .ZN(MRxD_Lb_1) );
  INV_X1 U28110 ( .A(1'b1), .ZN(MRxD_Lb_0) );
  INV_X1 U28112 ( .A(1'b1), .ZN(p_rxethmac1_LatchedByte_7) );
  INV_X1 U28114 ( .A(1'b1), .ZN(p_rxethmac1_LatchedByte_6) );
  INV_X1 U28116 ( .A(1'b1), .ZN(p_rxethmac1_LatchedByte_5) );
  INV_X1 U28118 ( .A(1'b1), .ZN(p_rxethmac1_LatchedByte_4) );
  INV_X1 U28120 ( .A(1'b1), .ZN(RxStateData_0) );
  INV_X1 U28122 ( .A(1'b1), .ZN(p_rxethmac1_n96) );
  INV_X1 U28124 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_0) );
  INV_X1 U28126 ( .A(1'b1), .ZN(p_rxethmac1_n97) );
  INV_X1 U28128 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_1) );
  INV_X1 U28130 ( .A(1'b1), .ZN(p_rxethmac1_n98) );
  INV_X1 U28132 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_2) );
  INV_X1 U28134 ( .A(1'b1), .ZN(p_rxethmac1_n99) );
  INV_X1 U28136 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_3) );
  INV_X1 U28138 ( .A(1'b1), .ZN(p_rxethmac1_n100) );
  INV_X1 U28140 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_4) );
  INV_X1 U28142 ( .A(1'b1), .ZN(p_rxethmac1_n101) );
  INV_X1 U28144 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_5) );
  INV_X1 U28146 ( .A(1'b1), .ZN(p_rxethmac1_n102) );
  INV_X1 U28148 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_6) );
  INV_X1 U28150 ( .A(1'b1), .ZN(p_rxethmac1_n103) );
  INV_X1 U28152 ( .A(1'b1), .ZN(p_rxethmac1_RxData_d_7) );
  INV_X1 U28154 ( .A(1'b0), .ZN(n33940) );
  INV_X1 U28156 ( .A(1'b0), .ZN(p_rxethmac1_GenerateRxStartFrm) );
  INV_X1 U28158 ( .A(1'b1), .ZN(p_rxethmac1_GenerateRxEndFrm) );
  INV_X1 U28160 ( .A(1'b0), .ZN(p_txethmac1_n154) );
  INV_X1 U28162 ( .A(1'b0), .ZN(p_txethmac1_n151) );
  INV_X1 U28164 ( .A(1'b0), .ZN(p_txethmac1_n156) );
  INV_X1 U28166 ( .A(1'b0), .ZN(p_txethmac1_n155) );
  INV_X1 U28168 ( .A(1'b0), .ZN(p_txethmac1_n150) );
  INV_X1 U28170 ( .A(1'b0), .ZN(p_txethmac1_n147) );
  INV_X1 U28172 ( .A(1'b0), .ZN(p_txethmac1_n148) );
  INV_X1 U28174 ( .A(1'b0), .ZN(p_txethmac1_n149) );
  INV_X1 U28176 ( .A(1'b1), .ZN(p_txethmac1_n153) );
  INV_X1 U28178 ( .A(1'b1), .ZN(p_txethmac1_n152) );
  INV_X1 U28180 ( .A(1'b0), .ZN(p_maccontrol1_n55) );
  INV_X1 U28182 ( .A(1'b1), .ZN(TxAbortIn) );
  INV_X1 U28184 ( .A(1'b1), .ZN(TxDoneIn) );
  INV_X1 U28186 ( .A(1'b0), .ZN(p_ethreg1_n686) );
  INV_X1 U28188 ( .A(1'b1), .ZN(p_ethreg1_SetTxCIrq_txclk) );
  INV_X1 U28190 ( .A(1'b1), .ZN(p_ethreg1_SetTxCIrq_sync2) );
  INV_X1 U28192 ( .A(1'b0), .ZN(p_ethreg1_N222) );
  INV_X1 U28194 ( .A(1'b1), .ZN(p_ethreg1_n685) );
  INV_X1 U28196 ( .A(1'b1), .ZN(p_ethreg1_SetRxCIrq_rxclk) );
  INV_X1 U28198 ( .A(1'b1), .ZN(p_ethreg1_SetRxCIrq_sync2) );
  INV_X1 U28200 ( .A(1'b0), .ZN(p_ethreg1_N228) );
  INV_X1 U28202 ( .A(1'b0), .ZN(p_ethreg1_n680) );
  INV_X1 U28204 ( .A(1'b1), .ZN(r_ScanStat) );
  INV_X1 U28206 ( .A(1'b0), .ZN(p_miim1_n152) );
  INV_X1 U28208 ( .A(1'b1), .ZN(r_RStat) );
  INV_X1 U28210 ( .A(1'b1), .ZN(p_miim1_RStat_q2) );
  INV_X1 U28212 ( .A(1'b1), .ZN(r_WCtrlData) );
  INV_X1 U28214 ( .A(1'b1), .ZN(p_miim1_WCtrlData_q2) );
  INV_X1 U28216 ( .A(1'b0), .ZN(p_miim1_n151) );
  INV_X1 U28218 ( .A(1'b1), .ZN(p_miim1_n150) );
  INV_X1 U28220 ( .A(1'b0), .ZN(p_miim1_n148) );
  INV_X1 U28222 ( .A(1'b0), .ZN(p_miim1_n155) );
  INV_X1 U28224 ( .A(1'b0), .ZN(p_miim1_n147) );
  INV_X1 U28226 ( .A(1'b0), .ZN(p_miim1_n146) );
  INV_X1 U28228 ( .A(1'b0), .ZN(p_miim1_n154) );
  INV_X1 U28230 ( .A(1'b0), .ZN(p_miim1_n145) );
  INV_X1 U28232 ( .A(1'b1), .ZN(p_miim1_n141) );
  INV_X1 U28234 ( .A(1'b0), .ZN(p_miim1_n139) );
  INV_X1 U28236 ( .A(1'b0), .ZN(p_miim1_n133) );
  INV_X1 U28238 ( .A(1'b0), .ZN(n124) );
  INV_X1 U28240 ( .A(1'b1), .ZN(WillSendControlFrame) );
  INV_X1 U28242 ( .A(1'b1), .ZN(md_padoe_o) );
  INV_X1 U28244 ( .A(1'b1), .ZN(md_pad_o) );
  INV_X1 U28246 ( .A(1'b1), .ZN(mdc_pad_o) );
  INV_X1 U28248 ( .A(1'b1), .ZN(mtxerr_pad_o) );
  INV_X1 U28250 ( .A(1'b1), .ZN(mtxen_pad_o) );
  INV_X1 U28252 ( .A(1'b1), .ZN(m_wb_stb_o) );
  INV_X1 U28254 ( .A(1'b1), .ZN(m_wb_cyc_o) );
  INV_X1 U28256 ( .A(1'b1), .ZN(m_wb_we_o) );
  INV_X1 U28258 ( .A(1'b1), .ZN(wb_err_o) );
  INV_X1 U28260 ( .A(1'b1), .ZN(wb_ack_o) );
  INV_X1 U28262 ( .A(1'b1), .ZN(mtxd_pad_o_3) );
  INV_X1 U28264 ( .A(1'b1), .ZN(mtxd_pad_o_2) );
  INV_X1 U28266 ( .A(1'b1), .ZN(mtxd_pad_o_1) );
  INV_X1 U28268 ( .A(1'b1), .ZN(mtxd_pad_o_0) );
  INV_X1 U28270 ( .A(1'b1), .ZN(m_wb_sel_o_3) );
  INV_X1 U28272 ( .A(1'b1), .ZN(m_wb_sel_o_2) );
  INV_X1 U28274 ( .A(1'b1), .ZN(m_wb_sel_o_1) );
  INV_X1 U28276 ( .A(1'b1), .ZN(m_wb_sel_o_0) );
  INV_X1 U28278 ( .A(1'b1), .ZN(m_wb_adr_o_31) );
  INV_X1 U28280 ( .A(1'b1), .ZN(m_wb_adr_o_30) );
  INV_X1 U28282 ( .A(1'b1), .ZN(m_wb_adr_o_29) );
  INV_X1 U28284 ( .A(1'b1), .ZN(m_wb_adr_o_28) );
  INV_X1 U28286 ( .A(1'b1), .ZN(m_wb_adr_o_27) );
  INV_X1 U28288 ( .A(1'b1), .ZN(m_wb_adr_o_26) );
  INV_X1 U28290 ( .A(1'b1), .ZN(m_wb_adr_o_25) );
  INV_X1 U28292 ( .A(1'b1), .ZN(m_wb_adr_o_24) );
  INV_X1 U28294 ( .A(1'b1), .ZN(m_wb_adr_o_23) );
  INV_X1 U28296 ( .A(1'b1), .ZN(m_wb_adr_o_22) );
  INV_X1 U28298 ( .A(1'b1), .ZN(m_wb_adr_o_21) );
  INV_X1 U28300 ( .A(1'b1), .ZN(m_wb_adr_o_20) );
  INV_X1 U28302 ( .A(1'b1), .ZN(m_wb_adr_o_19) );
  INV_X1 U28304 ( .A(1'b1), .ZN(m_wb_adr_o_18) );
  INV_X1 U28306 ( .A(1'b1), .ZN(m_wb_adr_o_17) );
  INV_X1 U28308 ( .A(1'b1), .ZN(m_wb_adr_o_16) );
  INV_X1 U28310 ( .A(1'b1), .ZN(m_wb_adr_o_15) );
  INV_X1 U28312 ( .A(1'b1), .ZN(m_wb_adr_o_14) );
  INV_X1 U28314 ( .A(1'b1), .ZN(m_wb_adr_o_13) );
  INV_X1 U28316 ( .A(1'b1), .ZN(m_wb_adr_o_12) );
  INV_X1 U28318 ( .A(1'b1), .ZN(m_wb_adr_o_11) );
  INV_X1 U28320 ( .A(1'b1), .ZN(m_wb_adr_o_10) );
  INV_X1 U28322 ( .A(1'b1), .ZN(m_wb_adr_o_9) );
  INV_X1 U28324 ( .A(1'b1), .ZN(m_wb_adr_o_8) );
  INV_X1 U28326 ( .A(1'b1), .ZN(m_wb_adr_o_7) );
  INV_X1 U28328 ( .A(1'b1), .ZN(m_wb_adr_o_6) );
  INV_X1 U28330 ( .A(1'b1), .ZN(m_wb_adr_o_5) );
  INV_X1 U28332 ( .A(1'b1), .ZN(m_wb_adr_o_4) );
  INV_X1 U28334 ( .A(1'b1), .ZN(m_wb_adr_o_3) );
  INV_X1 U28336 ( .A(1'b1), .ZN(m_wb_adr_o_2) );
  INV_X1 U28338 ( .A(1'b1), .ZN(m_wb_adr_o_1) );
  INV_X1 U28340 ( .A(1'b1), .ZN(m_wb_adr_o_0) );
  INV_X1 U28342 ( .A(n56254), .ZN(n23872) );
  INV_X1 U28343 ( .A(n23872), .ZN(temp_wb_dat_o_6) );
  INV_X1 U28344 ( .A(n56253), .ZN(n23874) );
  INV_X1 U28345 ( .A(n23874), .ZN(temp_wb_dat_o_5) );
  INV_X1 U28346 ( .A(n56252), .ZN(n23876) );
  INV_X1 U28347 ( .A(n23876), .ZN(temp_wb_dat_o_4) );
  INV_X1 U28348 ( .A(n56270), .ZN(n23878) );
  INV_X1 U28349 ( .A(n23878), .ZN(temp_wb_dat_o_31) );
  INV_X1 U28350 ( .A(n56269), .ZN(n23880) );
  INV_X1 U28351 ( .A(n23880), .ZN(temp_wb_dat_o_30) );
  INV_X1 U28352 ( .A(n56251), .ZN(n23882) );
  INV_X1 U28353 ( .A(n23882), .ZN(temp_wb_dat_o_3) );
  INV_X1 U28354 ( .A(n56268), .ZN(n23884) );
  INV_X1 U28355 ( .A(n23884), .ZN(temp_wb_dat_o_29) );
  INV_X1 U28356 ( .A(n56267), .ZN(n23886) );
  INV_X1 U28357 ( .A(n23886), .ZN(temp_wb_dat_o_28) );
  INV_X1 U28358 ( .A(n56266), .ZN(n23888) );
  INV_X1 U28359 ( .A(n23888), .ZN(temp_wb_dat_o_27) );
  INV_X1 U28360 ( .A(n56265), .ZN(n23890) );
  INV_X1 U28361 ( .A(n23890), .ZN(temp_wb_dat_o_26) );
  INV_X1 U28362 ( .A(n56264), .ZN(n23892) );
  INV_X1 U28363 ( .A(n23892), .ZN(temp_wb_dat_o_25) );
  INV_X1 U28364 ( .A(n56263), .ZN(n23894) );
  INV_X1 U28365 ( .A(n23894), .ZN(temp_wb_dat_o_24) );
  INV_X1 U28366 ( .A(n56262), .ZN(n23896) );
  INV_X1 U28367 ( .A(n23896), .ZN(temp_wb_dat_o_23) );
  INV_X1 U28368 ( .A(n56261), .ZN(n23898) );
  INV_X1 U28369 ( .A(n23898), .ZN(temp_wb_dat_o_22) );
  INV_X1 U28370 ( .A(n56260), .ZN(n23900) );
  INV_X1 U28371 ( .A(n23900), .ZN(temp_wb_dat_o_21) );
  INV_X1 U28372 ( .A(n56259), .ZN(n23902) );
  INV_X1 U28373 ( .A(n23902), .ZN(temp_wb_dat_o_20) );
  INV_X1 U28374 ( .A(n56250), .ZN(n23904) );
  INV_X1 U28375 ( .A(n23904), .ZN(temp_wb_dat_o_2) );
  INV_X1 U28376 ( .A(n56258), .ZN(n23906) );
  INV_X1 U28377 ( .A(n23906), .ZN(temp_wb_dat_o_19) );
  INV_X1 U28378 ( .A(n56257), .ZN(n23908) );
  INV_X1 U28379 ( .A(n23908), .ZN(temp_wb_dat_o_18) );
  INV_X1 U28380 ( .A(n56256), .ZN(n23910) );
  INV_X1 U28381 ( .A(n23910), .ZN(temp_wb_dat_o_17) );
  INV_X1 U28382 ( .A(n56255), .ZN(n23912) );
  INV_X1 U28383 ( .A(n23912), .ZN(temp_wb_dat_o_16) );
  INV_X1 U28384 ( .A(n56249), .ZN(n23914) );
  INV_X1 U28385 ( .A(n23914), .ZN(temp_wb_dat_o_1) );
  INV_X1 U28386 ( .A(n56248), .ZN(n23916) );
  INV_X1 U28387 ( .A(n23916), .ZN(temp_wb_dat_o_0) );
  INV_X1 U28388 ( .A(n64461), .ZN(n23918) );
  INV_X1 U28389 ( .A(n23918), .ZN(n34456) );
  INV_X1 U28390 ( .A(n32001), .ZN(n23920) );
  INV_X1 U28391 ( .A(n23920), .ZN(p_maccontrol1_transmitcontrol1_n279) );
  INV_X1 U28392 ( .A(n31388), .ZN(n23922) );
  INV_X1 U28393 ( .A(n23922), .ZN(p_miim1_shftrg_n140) );
  INV_X1 U28394 ( .A(n31377), .ZN(n23924) );
  INV_X1 U28395 ( .A(n23924), .ZN(p_miim1_shftrg_n141) );
  INV_X1 U28396 ( .A(n31365), .ZN(n23926) );
  INV_X1 U28397 ( .A(n23926), .ZN(p_miim1_shftrg_n142) );
  INV_X1 U28398 ( .A(n31354), .ZN(n23928) );
  INV_X1 U28399 ( .A(n23928), .ZN(p_miim1_shftrg_n143) );
  INV_X1 U28400 ( .A(n31339), .ZN(n23930) );
  INV_X1 U28401 ( .A(n23930), .ZN(p_miim1_shftrg_n144) );
  INV_X1 U28402 ( .A(n56246), .ZN(n23932) );
  INV_X1 U28403 ( .A(n23932), .ZN(n126) );
  INV_X1 U28404 ( .A(n56244), .ZN(n23934) );
  INV_X1 U28405 ( .A(n23934), .ZN(int_o) );
  INV_X1 U28406 ( .A(n64124), .ZN(n23936) );
  INV_X1 U28407 ( .A(n23936), .ZN(p_wishbone_tx_fifo_n1748) );
  INV_X1 U28408 ( .A(n64122), .ZN(n23938) );
  INV_X1 U28409 ( .A(n23938), .ZN(p_wishbone_tx_fifo_n1741) );
  INV_X1 U28410 ( .A(n56478), .ZN(n23940) );
  INV_X1 U28411 ( .A(n23940), .ZN(p_wishbone_n2472) );
  INV_X1 U28412 ( .A(n56396), .ZN(n23942) );
  INV_X1 U28413 ( .A(n23942), .ZN(p_wishbone_n2469) );
  INV_X1 U28414 ( .A(n56464), .ZN(n23944) );
  INV_X1 U28415 ( .A(n23944), .ZN(p_wishbone_n2467) );
  INV_X1 U28416 ( .A(n56460), .ZN(n23946) );
  INV_X1 U28417 ( .A(n23946), .ZN(p_wishbone_n2460) );
  INV_X1 U28418 ( .A(n56459), .ZN(n23948) );
  INV_X1 U28419 ( .A(n23948), .ZN(p_wishbone_n2458) );
  INV_X1 U28420 ( .A(n56397), .ZN(n23950) );
  INV_X1 U28421 ( .A(n23950), .ZN(p_wishbone_n2456) );
  INV_X1 U28422 ( .A(n56398), .ZN(n23952) );
  INV_X1 U28423 ( .A(n23952), .ZN(p_wishbone_n2455) );
  INV_X1 U28424 ( .A(n56399), .ZN(n23954) );
  INV_X1 U28425 ( .A(n23954), .ZN(p_wishbone_n2454) );
  INV_X1 U28426 ( .A(n56400), .ZN(n23956) );
  INV_X1 U28427 ( .A(n23956), .ZN(p_wishbone_n2453) );
  INV_X1 U28428 ( .A(n56401), .ZN(n23958) );
  INV_X1 U28429 ( .A(n23958), .ZN(p_wishbone_n2452) );
  INV_X1 U28430 ( .A(n56402), .ZN(n23960) );
  INV_X1 U28431 ( .A(n23960), .ZN(p_wishbone_n2451) );
  INV_X1 U28432 ( .A(n56403), .ZN(n23962) );
  INV_X1 U28433 ( .A(n23962), .ZN(p_wishbone_n2450) );
  INV_X1 U28434 ( .A(n56404), .ZN(n23964) );
  INV_X1 U28435 ( .A(n23964), .ZN(p_wishbone_n2449) );
  INV_X1 U28436 ( .A(n56405), .ZN(n23966) );
  INV_X1 U28437 ( .A(n23966), .ZN(p_wishbone_n2448) );
  INV_X1 U28438 ( .A(n56406), .ZN(n23968) );
  INV_X1 U28439 ( .A(n23968), .ZN(p_wishbone_n2447) );
  INV_X1 U28440 ( .A(n56407), .ZN(n23970) );
  INV_X1 U28441 ( .A(n23970), .ZN(p_wishbone_n2446) );
  INV_X1 U28442 ( .A(n56408), .ZN(n23972) );
  INV_X1 U28443 ( .A(n23972), .ZN(p_wishbone_n2445) );
  INV_X1 U28444 ( .A(n56409), .ZN(n23974) );
  INV_X1 U28445 ( .A(n23974), .ZN(p_wishbone_n2444) );
  INV_X1 U28446 ( .A(n56410), .ZN(n23976) );
  INV_X1 U28447 ( .A(n23976), .ZN(p_wishbone_n2443) );
  INV_X1 U28448 ( .A(n56411), .ZN(n23978) );
  INV_X1 U28449 ( .A(n23978), .ZN(p_wishbone_n2442) );
  INV_X1 U28450 ( .A(n56394), .ZN(n23980) );
  INV_X1 U28451 ( .A(n23980), .ZN(p_wishbone_n2441) );
  INV_X1 U28452 ( .A(n56412), .ZN(n23982) );
  INV_X1 U28453 ( .A(n23982), .ZN(p_wishbone_n2440) );
  INV_X1 U28454 ( .A(n56413), .ZN(n23984) );
  INV_X1 U28455 ( .A(n23984), .ZN(p_wishbone_n2439) );
  INV_X1 U28456 ( .A(n56414), .ZN(n23986) );
  INV_X1 U28457 ( .A(n23986), .ZN(p_wishbone_n2438) );
  INV_X1 U28458 ( .A(n56380), .ZN(n23988) );
  INV_X1 U28459 ( .A(n23988), .ZN(p_wishbone_n2437) );
  INV_X1 U28460 ( .A(n56415), .ZN(n23990) );
  INV_X1 U28461 ( .A(n23990), .ZN(p_wishbone_n2436) );
  INV_X1 U28462 ( .A(n56470), .ZN(n23992) );
  INV_X1 U28463 ( .A(n23992), .ZN(p_wishbone_n2435) );
  INV_X1 U28464 ( .A(n56416), .ZN(n23994) );
  INV_X1 U28465 ( .A(n23994), .ZN(p_wishbone_n2434) );
  INV_X1 U28466 ( .A(n56417), .ZN(n23996) );
  INV_X1 U28467 ( .A(n23996), .ZN(p_wishbone_n2433) );
  INV_X1 U28468 ( .A(n56418), .ZN(n23998) );
  INV_X1 U28469 ( .A(n23998), .ZN(p_wishbone_n2432) );
  INV_X1 U28470 ( .A(n56419), .ZN(n24000) );
  INV_X1 U28471 ( .A(n24000), .ZN(p_wishbone_n2431) );
  INV_X1 U28472 ( .A(n56420), .ZN(n24002) );
  INV_X1 U28473 ( .A(n24002), .ZN(p_wishbone_n2430) );
  INV_X1 U28474 ( .A(n56421), .ZN(n24004) );
  INV_X1 U28475 ( .A(n24004), .ZN(p_wishbone_n2429) );
  INV_X1 U28476 ( .A(n56438), .ZN(n24006) );
  INV_X1 U28477 ( .A(n24006), .ZN(p_wishbone_n2426) );
  INV_X1 U28478 ( .A(n56427), .ZN(n24008) );
  INV_X1 U28479 ( .A(n24008), .ZN(p_wishbone_n2423) );
  INV_X1 U28480 ( .A(n56426), .ZN(n24010) );
  INV_X1 U28481 ( .A(n24010), .ZN(p_wishbone_n2422) );
  INV_X1 U28482 ( .A(n56425), .ZN(n24012) );
  INV_X1 U28483 ( .A(n24012), .ZN(p_wishbone_n2421) );
  INV_X1 U28484 ( .A(n56424), .ZN(n24014) );
  INV_X1 U28485 ( .A(n24014), .ZN(p_wishbone_n2420) );
  INV_X1 U28486 ( .A(n56423), .ZN(n24016) );
  INV_X1 U28487 ( .A(n24016), .ZN(p_wishbone_n2419) );
  INV_X1 U28488 ( .A(n56422), .ZN(n24018) );
  INV_X1 U28489 ( .A(n24018), .ZN(p_wishbone_n2418) );
  INV_X1 U28490 ( .A(n56430), .ZN(n24020) );
  INV_X1 U28491 ( .A(n24020), .ZN(p_wishbone_n2411) );
  INV_X1 U28492 ( .A(n56437), .ZN(n24022) );
  INV_X1 U28493 ( .A(n24022), .ZN(p_wishbone_n2409) );
  INV_X1 U28494 ( .A(n56436), .ZN(n24024) );
  INV_X1 U28495 ( .A(n24024), .ZN(p_wishbone_n2408) );
  INV_X1 U28496 ( .A(n56462), .ZN(n24026) );
  INV_X1 U28497 ( .A(n24026), .ZN(p_wishbone_n2350) );
  INV_X1 U28498 ( .A(n56372), .ZN(n24028) );
  INV_X1 U28499 ( .A(n24028), .ZN(p_wishbone_n2334) );
  INV_X1 U28500 ( .A(n56440), .ZN(n24030) );
  INV_X1 U28501 ( .A(n24030), .ZN(p_wishbone_n2332) );
  INV_X1 U28502 ( .A(n56457), .ZN(n24032) );
  INV_X1 U28503 ( .A(n24032), .ZN(p_wishbone_n2316) );
  INV_X1 U28504 ( .A(n56456), .ZN(n24034) );
  INV_X1 U28505 ( .A(n24034), .ZN(p_wishbone_n2315) );
  INV_X1 U28506 ( .A(n56455), .ZN(n24036) );
  INV_X1 U28507 ( .A(n24036), .ZN(p_wishbone_n2314) );
  INV_X1 U28508 ( .A(n56454), .ZN(n24038) );
  INV_X1 U28509 ( .A(n24038), .ZN(p_wishbone_n2313) );
  INV_X1 U28510 ( .A(n56453), .ZN(n24040) );
  INV_X1 U28511 ( .A(n24040), .ZN(p_wishbone_n2312) );
  INV_X1 U28512 ( .A(n56452), .ZN(n24042) );
  INV_X1 U28513 ( .A(n24042), .ZN(p_wishbone_n2311) );
  INV_X1 U28514 ( .A(n56451), .ZN(n24044) );
  INV_X1 U28515 ( .A(n24044), .ZN(p_wishbone_n2310) );
  INV_X1 U28516 ( .A(n56450), .ZN(n24046) );
  INV_X1 U28517 ( .A(n24046), .ZN(p_wishbone_n2309) );
  INV_X1 U28518 ( .A(n56449), .ZN(n24048) );
  INV_X1 U28519 ( .A(n24048), .ZN(p_wishbone_n2308) );
  INV_X1 U28520 ( .A(n56448), .ZN(n24050) );
  INV_X1 U28521 ( .A(n24050), .ZN(p_wishbone_n2307) );
  INV_X1 U28522 ( .A(n56447), .ZN(n24052) );
  INV_X1 U28523 ( .A(n24052), .ZN(p_wishbone_n2306) );
  INV_X1 U28524 ( .A(n56446), .ZN(n24054) );
  INV_X1 U28525 ( .A(n24054), .ZN(p_wishbone_n2305) );
  INV_X1 U28526 ( .A(n56445), .ZN(n24056) );
  INV_X1 U28527 ( .A(n24056), .ZN(p_wishbone_n2304) );
  INV_X1 U28528 ( .A(n56444), .ZN(n24058) );
  INV_X1 U28529 ( .A(n24058), .ZN(p_wishbone_n2303) );
  INV_X1 U28530 ( .A(n56443), .ZN(n24060) );
  INV_X1 U28531 ( .A(n24060), .ZN(p_wishbone_n2302) );
  INV_X1 U28532 ( .A(n56468), .ZN(n24062) );
  INV_X1 U28533 ( .A(n24062), .ZN(p_wishbone_n2297) );
  INV_X1 U28534 ( .A(n56377), .ZN(n24064) );
  INV_X1 U28535 ( .A(n24064), .ZN(p_wishbone_n2292) );
  INV_X1 U28536 ( .A(n56376), .ZN(n24066) );
  INV_X1 U28537 ( .A(n24066), .ZN(p_wishbone_n2253) );
  INV_X1 U28538 ( .A(n56375), .ZN(n24068) );
  INV_X1 U28539 ( .A(n24068), .ZN(p_wishbone_n2252) );
  INV_X1 U28540 ( .A(n56374), .ZN(n24070) );
  INV_X1 U28541 ( .A(n24070), .ZN(p_wishbone_n2251) );
  INV_X1 U28542 ( .A(n56373), .ZN(n24072) );
  INV_X1 U28543 ( .A(n24072), .ZN(p_wishbone_n2250) );
  INV_X1 U28544 ( .A(n56442), .ZN(n24074) );
  INV_X1 U28545 ( .A(n24074), .ZN(p_wishbone_n2248) );
  INV_X1 U28546 ( .A(n56393), .ZN(n24076) );
  INV_X1 U28547 ( .A(n24076), .ZN(p_wishbone_n2240) );
  INV_X1 U28548 ( .A(n56386), .ZN(n24078) );
  INV_X1 U28549 ( .A(n24078), .ZN(p_wishbone_n2239) );
  INV_X1 U28550 ( .A(n56392), .ZN(n24080) );
  INV_X1 U28551 ( .A(n24080), .ZN(p_wishbone_n2238) );
  INV_X1 U28552 ( .A(n56391), .ZN(n24082) );
  INV_X1 U28553 ( .A(n24082), .ZN(p_wishbone_n2237) );
  INV_X1 U28554 ( .A(n56390), .ZN(n24084) );
  INV_X1 U28555 ( .A(n24084), .ZN(p_wishbone_n2236) );
  INV_X1 U28556 ( .A(n56389), .ZN(n24086) );
  INV_X1 U28557 ( .A(n24086), .ZN(p_wishbone_n2235) );
  INV_X1 U28558 ( .A(n56388), .ZN(n24088) );
  INV_X1 U28559 ( .A(n24088), .ZN(p_wishbone_n2234) );
  INV_X1 U28560 ( .A(n56387), .ZN(n24090) );
  INV_X1 U28561 ( .A(n24090), .ZN(p_wishbone_n2233) );
  INV_X1 U28562 ( .A(n56381), .ZN(n24092) );
  INV_X1 U28563 ( .A(n24092), .ZN(p_wishbone_n2231) );
  INV_X1 U28564 ( .A(n56370), .ZN(n24094) );
  INV_X1 U28565 ( .A(n24094), .ZN(p_wishbone_n2229) );
  INV_X1 U28566 ( .A(n56369), .ZN(n24096) );
  INV_X1 U28567 ( .A(n24096), .ZN(p_wishbone_n2228) );
  INV_X1 U28568 ( .A(n56368), .ZN(n24098) );
  INV_X1 U28569 ( .A(n24098), .ZN(p_wishbone_n2227) );
  INV_X1 U28570 ( .A(n56367), .ZN(n24100) );
  INV_X1 U28571 ( .A(n24100), .ZN(p_wishbone_n2226) );
  INV_X1 U28572 ( .A(n56366), .ZN(n24102) );
  INV_X1 U28573 ( .A(n24102), .ZN(p_wishbone_n2225) );
  INV_X1 U28574 ( .A(n56365), .ZN(n24104) );
  INV_X1 U28575 ( .A(n24104), .ZN(p_wishbone_n2224) );
  INV_X1 U28576 ( .A(n56364), .ZN(n24106) );
  INV_X1 U28577 ( .A(n24106), .ZN(p_wishbone_n2223) );
  INV_X1 U28578 ( .A(n56363), .ZN(n24108) );
  INV_X1 U28579 ( .A(n24108), .ZN(p_wishbone_n2222) );
  INV_X1 U28580 ( .A(n56362), .ZN(n24110) );
  INV_X1 U28581 ( .A(n24110), .ZN(p_wishbone_n2221) );
  INV_X1 U28582 ( .A(n56361), .ZN(n24112) );
  INV_X1 U28583 ( .A(n24112), .ZN(p_wishbone_n2220) );
  INV_X1 U28584 ( .A(n56360), .ZN(n24114) );
  INV_X1 U28585 ( .A(n24114), .ZN(p_wishbone_n2219) );
  INV_X1 U28586 ( .A(n56359), .ZN(n24116) );
  INV_X1 U28587 ( .A(n24116), .ZN(p_wishbone_n2218) );
  INV_X1 U28588 ( .A(n56358), .ZN(n24118) );
  INV_X1 U28589 ( .A(n24118), .ZN(p_wishbone_n2217) );
  INV_X1 U28590 ( .A(n56357), .ZN(n24120) );
  INV_X1 U28591 ( .A(n24120), .ZN(p_wishbone_n2216) );
  INV_X1 U28592 ( .A(n56356), .ZN(n24122) );
  INV_X1 U28593 ( .A(n24122), .ZN(p_wishbone_n2215) );
  INV_X1 U28594 ( .A(n56355), .ZN(n24124) );
  INV_X1 U28595 ( .A(n24124), .ZN(p_wishbone_n2214) );
  INV_X1 U28596 ( .A(n56354), .ZN(n24126) );
  INV_X1 U28597 ( .A(n24126), .ZN(p_wishbone_n2213) );
  INV_X1 U28598 ( .A(n56353), .ZN(n24128) );
  INV_X1 U28599 ( .A(n24128), .ZN(p_wishbone_n2212) );
  INV_X1 U28600 ( .A(n56352), .ZN(n24130) );
  INV_X1 U28601 ( .A(n24130), .ZN(p_wishbone_n2211) );
  INV_X1 U28602 ( .A(n56351), .ZN(n24132) );
  INV_X1 U28603 ( .A(n24132), .ZN(p_wishbone_n2210) );
  INV_X1 U28604 ( .A(n56350), .ZN(n24134) );
  INV_X1 U28605 ( .A(n24134), .ZN(p_wishbone_n2209) );
  INV_X1 U28606 ( .A(n56349), .ZN(n24136) );
  INV_X1 U28607 ( .A(n24136), .ZN(p_wishbone_n2208) );
  INV_X1 U28608 ( .A(n56348), .ZN(n24138) );
  INV_X1 U28609 ( .A(n24138), .ZN(p_wishbone_n2207) );
  INV_X1 U28610 ( .A(n56347), .ZN(n24140) );
  INV_X1 U28611 ( .A(n24140), .ZN(p_wishbone_n2206) );
  INV_X1 U28612 ( .A(n56346), .ZN(n24142) );
  INV_X1 U28613 ( .A(n24142), .ZN(p_wishbone_n2205) );
  INV_X1 U28614 ( .A(n56345), .ZN(n24144) );
  INV_X1 U28615 ( .A(n24144), .ZN(p_wishbone_n2204) );
  INV_X1 U28616 ( .A(n56344), .ZN(n24146) );
  INV_X1 U28617 ( .A(n24146), .ZN(p_wishbone_n2203) );
  INV_X1 U28618 ( .A(n56343), .ZN(n24148) );
  INV_X1 U28619 ( .A(n24148), .ZN(p_wishbone_n2202) );
  INV_X1 U28620 ( .A(n56342), .ZN(n24150) );
  INV_X1 U28621 ( .A(n24150), .ZN(p_wishbone_n2201) );
  INV_X1 U28622 ( .A(n56371), .ZN(n24152) );
  INV_X1 U28623 ( .A(n24152), .ZN(p_wishbone_n2200) );
  INV_X1 U28624 ( .A(n56340), .ZN(n24154) );
  INV_X1 U28625 ( .A(n24154), .ZN(p_wishbone_n2199) );
  INV_X1 U28626 ( .A(n56339), .ZN(n24156) );
  INV_X1 U28627 ( .A(n24156), .ZN(p_wishbone_n2198) );
  INV_X1 U28628 ( .A(n56338), .ZN(n24158) );
  INV_X1 U28629 ( .A(n24158), .ZN(p_wishbone_n2197) );
  INV_X1 U28630 ( .A(n56337), .ZN(n24160) );
  INV_X1 U28631 ( .A(n24160), .ZN(p_wishbone_n2196) );
  INV_X1 U28632 ( .A(n56336), .ZN(n24162) );
  INV_X1 U28633 ( .A(n24162), .ZN(p_wishbone_n2195) );
  INV_X1 U28634 ( .A(n56335), .ZN(n24164) );
  INV_X1 U28635 ( .A(n24164), .ZN(p_wishbone_n2194) );
  INV_X1 U28636 ( .A(n56334), .ZN(n24166) );
  INV_X1 U28637 ( .A(n24166), .ZN(p_wishbone_n2193) );
  INV_X1 U28638 ( .A(n56333), .ZN(n24168) );
  INV_X1 U28639 ( .A(n24168), .ZN(p_wishbone_n2192) );
  INV_X1 U28640 ( .A(n56332), .ZN(n24170) );
  INV_X1 U28641 ( .A(n24170), .ZN(p_wishbone_n2191) );
  INV_X1 U28642 ( .A(n56331), .ZN(n24172) );
  INV_X1 U28643 ( .A(n24172), .ZN(p_wishbone_n2190) );
  INV_X1 U28644 ( .A(n56330), .ZN(n24174) );
  INV_X1 U28645 ( .A(n24174), .ZN(p_wishbone_n2189) );
  INV_X1 U28646 ( .A(n56329), .ZN(n24176) );
  INV_X1 U28647 ( .A(n24176), .ZN(p_wishbone_n2188) );
  INV_X1 U28648 ( .A(n56328), .ZN(n24178) );
  INV_X1 U28649 ( .A(n24178), .ZN(p_wishbone_n2187) );
  INV_X1 U28650 ( .A(n56327), .ZN(n24180) );
  INV_X1 U28651 ( .A(n24180), .ZN(p_wishbone_n2186) );
  INV_X1 U28652 ( .A(n56326), .ZN(n24182) );
  INV_X1 U28653 ( .A(n24182), .ZN(p_wishbone_n2185) );
  INV_X1 U28654 ( .A(n56325), .ZN(n24184) );
  INV_X1 U28655 ( .A(n24184), .ZN(p_wishbone_n2184) );
  INV_X1 U28656 ( .A(n56324), .ZN(n24186) );
  INV_X1 U28657 ( .A(n24186), .ZN(p_wishbone_n2183) );
  INV_X1 U28658 ( .A(n56323), .ZN(n24188) );
  INV_X1 U28659 ( .A(n24188), .ZN(p_wishbone_n2182) );
  INV_X1 U28660 ( .A(n56322), .ZN(n24190) );
  INV_X1 U28661 ( .A(n24190), .ZN(p_wishbone_n2181) );
  INV_X1 U28662 ( .A(n56321), .ZN(n24192) );
  INV_X1 U28663 ( .A(n24192), .ZN(p_wishbone_n2180) );
  INV_X1 U28664 ( .A(n56320), .ZN(n24194) );
  INV_X1 U28665 ( .A(n24194), .ZN(p_wishbone_n2179) );
  INV_X1 U28666 ( .A(n56319), .ZN(n24196) );
  INV_X1 U28667 ( .A(n24196), .ZN(p_wishbone_n2178) );
  INV_X1 U28668 ( .A(n56318), .ZN(n24198) );
  INV_X1 U28669 ( .A(n24198), .ZN(p_wishbone_n2177) );
  INV_X1 U28670 ( .A(n56317), .ZN(n24200) );
  INV_X1 U28671 ( .A(n24200), .ZN(p_wishbone_n2176) );
  INV_X1 U28672 ( .A(n56316), .ZN(n24202) );
  INV_X1 U28673 ( .A(n24202), .ZN(p_wishbone_n2175) );
  INV_X1 U28674 ( .A(n56315), .ZN(n24204) );
  INV_X1 U28675 ( .A(n24204), .ZN(p_wishbone_n2174) );
  INV_X1 U28676 ( .A(n56314), .ZN(n24206) );
  INV_X1 U28677 ( .A(n24206), .ZN(p_wishbone_n2173) );
  INV_X1 U28678 ( .A(n56313), .ZN(n24208) );
  INV_X1 U28679 ( .A(n24208), .ZN(p_wishbone_n2172) );
  INV_X1 U28680 ( .A(n56312), .ZN(n24210) );
  INV_X1 U28681 ( .A(n24210), .ZN(p_wishbone_n2171) );
  INV_X1 U28682 ( .A(n56341), .ZN(n24212) );
  INV_X1 U28683 ( .A(n24212), .ZN(p_wishbone_n2170) );
  INV_X1 U28684 ( .A(n56311), .ZN(n24214) );
  INV_X1 U28685 ( .A(n24214), .ZN(p_wishbone_n2142) );
  INV_X1 U28686 ( .A(n64121), .ZN(n24216) );
  INV_X1 U28687 ( .A(n24216), .ZN(p_wishbone_bd_ram_n25984) );
  INV_X1 U28688 ( .A(n64120), .ZN(n24218) );
  INV_X1 U28689 ( .A(n24218), .ZN(p_wishbone_bd_ram_n25983) );
  INV_X1 U28690 ( .A(n64119), .ZN(n24220) );
  INV_X1 U28691 ( .A(n24220), .ZN(p_wishbone_bd_ram_n25982) );
  INV_X1 U28692 ( .A(n64118), .ZN(n24222) );
  INV_X1 U28693 ( .A(n24222), .ZN(p_wishbone_bd_ram_n25981) );
  INV_X1 U28694 ( .A(n64117), .ZN(n24224) );
  INV_X1 U28695 ( .A(n24224), .ZN(p_wishbone_bd_ram_n25980) );
  INV_X1 U28696 ( .A(n64116), .ZN(n24226) );
  INV_X1 U28697 ( .A(n24226), .ZN(p_wishbone_bd_ram_n25979) );
  INV_X1 U28698 ( .A(n64115), .ZN(n24228) );
  INV_X1 U28699 ( .A(n24228), .ZN(p_wishbone_bd_ram_n25978) );
  INV_X1 U28700 ( .A(n64114), .ZN(n24230) );
  INV_X1 U28701 ( .A(n24230), .ZN(p_wishbone_bd_ram_n25977) );
  INV_X1 U28702 ( .A(n64113), .ZN(n24232) );
  INV_X1 U28703 ( .A(n24232), .ZN(p_wishbone_bd_ram_n25976) );
  INV_X1 U28704 ( .A(n64112), .ZN(n24234) );
  INV_X1 U28705 ( .A(n24234), .ZN(p_wishbone_bd_ram_n25975) );
  INV_X1 U28706 ( .A(n64111), .ZN(n24236) );
  INV_X1 U28707 ( .A(n24236), .ZN(p_wishbone_bd_ram_n25974) );
  INV_X1 U28708 ( .A(n64110), .ZN(n24238) );
  INV_X1 U28709 ( .A(n24238), .ZN(p_wishbone_bd_ram_n25973) );
  INV_X1 U28710 ( .A(n64109), .ZN(n24240) );
  INV_X1 U28711 ( .A(n24240), .ZN(p_wishbone_bd_ram_n25972) );
  INV_X1 U28712 ( .A(n64108), .ZN(n24242) );
  INV_X1 U28713 ( .A(n24242), .ZN(p_wishbone_bd_ram_n25971) );
  INV_X1 U28714 ( .A(n64107), .ZN(n24244) );
  INV_X1 U28715 ( .A(n24244), .ZN(p_wishbone_bd_ram_n25970) );
  INV_X1 U28716 ( .A(n64106), .ZN(n24246) );
  INV_X1 U28717 ( .A(n24246), .ZN(p_wishbone_bd_ram_n25969) );
  INV_X1 U28718 ( .A(n64105), .ZN(n24248) );
  INV_X1 U28719 ( .A(n24248), .ZN(p_wishbone_bd_ram_n25968) );
  INV_X1 U28720 ( .A(n64104), .ZN(n24250) );
  INV_X1 U28721 ( .A(n24250), .ZN(p_wishbone_bd_ram_n25967) );
  INV_X1 U28722 ( .A(n64103), .ZN(n24252) );
  INV_X1 U28723 ( .A(n24252), .ZN(p_wishbone_bd_ram_n25966) );
  INV_X1 U28724 ( .A(n64102), .ZN(n24254) );
  INV_X1 U28725 ( .A(n24254), .ZN(p_wishbone_bd_ram_n25965) );
  INV_X1 U28726 ( .A(n64101), .ZN(n24256) );
  INV_X1 U28727 ( .A(n24256), .ZN(p_wishbone_bd_ram_n25964) );
  INV_X1 U28728 ( .A(n64100), .ZN(n24258) );
  INV_X1 U28729 ( .A(n24258), .ZN(p_wishbone_bd_ram_n25963) );
  INV_X1 U28730 ( .A(n64099), .ZN(n24260) );
  INV_X1 U28731 ( .A(n24260), .ZN(p_wishbone_bd_ram_n25962) );
  INV_X1 U28732 ( .A(n64098), .ZN(n24262) );
  INV_X1 U28733 ( .A(n24262), .ZN(p_wishbone_bd_ram_n25961) );
  INV_X1 U28734 ( .A(n64097), .ZN(n24264) );
  INV_X1 U28735 ( .A(n24264), .ZN(p_wishbone_bd_ram_n25960) );
  INV_X1 U28736 ( .A(n64096), .ZN(n24266) );
  INV_X1 U28737 ( .A(n24266), .ZN(p_wishbone_bd_ram_n25959) );
  INV_X1 U28738 ( .A(n64095), .ZN(n24268) );
  INV_X1 U28739 ( .A(n24268), .ZN(p_wishbone_bd_ram_n25958) );
  INV_X1 U28740 ( .A(n64094), .ZN(n24270) );
  INV_X1 U28741 ( .A(n24270), .ZN(p_wishbone_bd_ram_n25957) );
  INV_X1 U28742 ( .A(n64093), .ZN(n24272) );
  INV_X1 U28743 ( .A(n24272), .ZN(p_wishbone_bd_ram_n25956) );
  INV_X1 U28744 ( .A(n64092), .ZN(n24274) );
  INV_X1 U28745 ( .A(n24274), .ZN(p_wishbone_bd_ram_n25955) );
  INV_X1 U28746 ( .A(n64091), .ZN(n24276) );
  INV_X1 U28747 ( .A(n24276), .ZN(p_wishbone_bd_ram_n25954) );
  INV_X1 U28748 ( .A(n64090), .ZN(n24278) );
  INV_X1 U28749 ( .A(n24278), .ZN(p_wishbone_bd_ram_n25953) );
  INV_X1 U28750 ( .A(n64089), .ZN(n24280) );
  INV_X1 U28751 ( .A(n24280), .ZN(p_wishbone_bd_ram_n25952) );
  INV_X1 U28752 ( .A(n64088), .ZN(n24282) );
  INV_X1 U28753 ( .A(n24282), .ZN(p_wishbone_bd_ram_n25951) );
  INV_X1 U28754 ( .A(n64087), .ZN(n24284) );
  INV_X1 U28755 ( .A(n24284), .ZN(p_wishbone_bd_ram_n25950) );
  INV_X1 U28756 ( .A(n64086), .ZN(n24286) );
  INV_X1 U28757 ( .A(n24286), .ZN(p_wishbone_bd_ram_n25949) );
  INV_X1 U28758 ( .A(n64085), .ZN(n24288) );
  INV_X1 U28759 ( .A(n24288), .ZN(p_wishbone_bd_ram_n25948) );
  INV_X1 U28760 ( .A(n64084), .ZN(n24290) );
  INV_X1 U28761 ( .A(n24290), .ZN(p_wishbone_bd_ram_n25947) );
  INV_X1 U28762 ( .A(n64083), .ZN(n24292) );
  INV_X1 U28763 ( .A(n24292), .ZN(p_wishbone_bd_ram_n25946) );
  INV_X1 U28764 ( .A(n64082), .ZN(n24294) );
  INV_X1 U28765 ( .A(n24294), .ZN(p_wishbone_bd_ram_n25945) );
  INV_X1 U28766 ( .A(n64081), .ZN(n24296) );
  INV_X1 U28767 ( .A(n24296), .ZN(p_wishbone_bd_ram_n25944) );
  INV_X1 U28768 ( .A(n64080), .ZN(n24298) );
  INV_X1 U28769 ( .A(n24298), .ZN(p_wishbone_bd_ram_n25943) );
  INV_X1 U28770 ( .A(n64079), .ZN(n24300) );
  INV_X1 U28771 ( .A(n24300), .ZN(p_wishbone_bd_ram_n25942) );
  INV_X1 U28772 ( .A(n64078), .ZN(n24302) );
  INV_X1 U28773 ( .A(n24302), .ZN(p_wishbone_bd_ram_n25941) );
  INV_X1 U28774 ( .A(n64077), .ZN(n24304) );
  INV_X1 U28775 ( .A(n24304), .ZN(p_wishbone_bd_ram_n25940) );
  INV_X1 U28776 ( .A(n64076), .ZN(n24306) );
  INV_X1 U28777 ( .A(n24306), .ZN(p_wishbone_bd_ram_n25939) );
  INV_X1 U28778 ( .A(n64075), .ZN(n24308) );
  INV_X1 U28779 ( .A(n24308), .ZN(p_wishbone_bd_ram_n25938) );
  INV_X1 U28780 ( .A(n64074), .ZN(n24310) );
  INV_X1 U28781 ( .A(n24310), .ZN(p_wishbone_bd_ram_n25937) );
  INV_X1 U28782 ( .A(n64073), .ZN(n24312) );
  INV_X1 U28783 ( .A(n24312), .ZN(p_wishbone_bd_ram_n25936) );
  INV_X1 U28784 ( .A(n64072), .ZN(n24314) );
  INV_X1 U28785 ( .A(n24314), .ZN(p_wishbone_bd_ram_n25935) );
  INV_X1 U28786 ( .A(n64071), .ZN(n24316) );
  INV_X1 U28787 ( .A(n24316), .ZN(p_wishbone_bd_ram_n25934) );
  INV_X1 U28788 ( .A(n64070), .ZN(n24318) );
  INV_X1 U28789 ( .A(n24318), .ZN(p_wishbone_bd_ram_n25933) );
  INV_X1 U28790 ( .A(n64069), .ZN(n24320) );
  INV_X1 U28791 ( .A(n24320), .ZN(p_wishbone_bd_ram_n25932) );
  INV_X1 U28792 ( .A(n64068), .ZN(n24322) );
  INV_X1 U28793 ( .A(n24322), .ZN(p_wishbone_bd_ram_n25931) );
  INV_X1 U28794 ( .A(n64067), .ZN(n24324) );
  INV_X1 U28795 ( .A(n24324), .ZN(p_wishbone_bd_ram_n25930) );
  INV_X1 U28796 ( .A(n64066), .ZN(n24326) );
  INV_X1 U28797 ( .A(n24326), .ZN(p_wishbone_bd_ram_n25929) );
  INV_X1 U28798 ( .A(n64065), .ZN(n24328) );
  INV_X1 U28799 ( .A(n24328), .ZN(p_wishbone_bd_ram_n25928) );
  INV_X1 U28800 ( .A(n64064), .ZN(n24330) );
  INV_X1 U28801 ( .A(n24330), .ZN(p_wishbone_bd_ram_n25927) );
  INV_X1 U28802 ( .A(n64063), .ZN(n24332) );
  INV_X1 U28803 ( .A(n24332), .ZN(p_wishbone_bd_ram_n25926) );
  INV_X1 U28804 ( .A(n64062), .ZN(n24334) );
  INV_X1 U28805 ( .A(n24334), .ZN(p_wishbone_bd_ram_n25925) );
  INV_X1 U28806 ( .A(n64061), .ZN(n24336) );
  INV_X1 U28807 ( .A(n24336), .ZN(p_wishbone_bd_ram_n25924) );
  INV_X1 U28808 ( .A(n64060), .ZN(n24338) );
  INV_X1 U28809 ( .A(n24338), .ZN(p_wishbone_bd_ram_n25923) );
  INV_X1 U28810 ( .A(n64059), .ZN(n24340) );
  INV_X1 U28811 ( .A(n24340), .ZN(p_wishbone_bd_ram_n25922) );
  INV_X1 U28812 ( .A(n64058), .ZN(n24342) );
  INV_X1 U28813 ( .A(n24342), .ZN(p_wishbone_bd_ram_n25921) );
  INV_X1 U28814 ( .A(n64057), .ZN(n24344) );
  INV_X1 U28815 ( .A(n24344), .ZN(p_wishbone_bd_ram_n25920) );
  INV_X1 U28816 ( .A(n64056), .ZN(n24346) );
  INV_X1 U28817 ( .A(n24346), .ZN(p_wishbone_bd_ram_n25919) );
  INV_X1 U28818 ( .A(n64055), .ZN(n24348) );
  INV_X1 U28819 ( .A(n24348), .ZN(p_wishbone_bd_ram_n25918) );
  INV_X1 U28820 ( .A(n64054), .ZN(n24350) );
  INV_X1 U28821 ( .A(n24350), .ZN(p_wishbone_bd_ram_n25917) );
  INV_X1 U28822 ( .A(n64053), .ZN(n24352) );
  INV_X1 U28823 ( .A(n24352), .ZN(p_wishbone_bd_ram_n25916) );
  INV_X1 U28824 ( .A(n64052), .ZN(n24354) );
  INV_X1 U28825 ( .A(n24354), .ZN(p_wishbone_bd_ram_n25915) );
  INV_X1 U28826 ( .A(n64051), .ZN(n24356) );
  INV_X1 U28827 ( .A(n24356), .ZN(p_wishbone_bd_ram_n25914) );
  INV_X1 U28828 ( .A(n64050), .ZN(n24358) );
  INV_X1 U28829 ( .A(n24358), .ZN(p_wishbone_bd_ram_n25913) );
  INV_X1 U28830 ( .A(n64049), .ZN(n24360) );
  INV_X1 U28831 ( .A(n24360), .ZN(p_wishbone_bd_ram_n25912) );
  INV_X1 U28832 ( .A(n64048), .ZN(n24362) );
  INV_X1 U28833 ( .A(n24362), .ZN(p_wishbone_bd_ram_n25911) );
  INV_X1 U28834 ( .A(n64047), .ZN(n24364) );
  INV_X1 U28835 ( .A(n24364), .ZN(p_wishbone_bd_ram_n25910) );
  INV_X1 U28836 ( .A(n64046), .ZN(n24366) );
  INV_X1 U28837 ( .A(n24366), .ZN(p_wishbone_bd_ram_n25909) );
  INV_X1 U28838 ( .A(n64045), .ZN(n24368) );
  INV_X1 U28839 ( .A(n24368), .ZN(p_wishbone_bd_ram_n25908) );
  INV_X1 U28840 ( .A(n64044), .ZN(n24370) );
  INV_X1 U28841 ( .A(n24370), .ZN(p_wishbone_bd_ram_n25907) );
  INV_X1 U28842 ( .A(n64043), .ZN(n24372) );
  INV_X1 U28843 ( .A(n24372), .ZN(p_wishbone_bd_ram_n25906) );
  INV_X1 U28844 ( .A(n64042), .ZN(n24374) );
  INV_X1 U28845 ( .A(n24374), .ZN(p_wishbone_bd_ram_n25905) );
  INV_X1 U28846 ( .A(n64041), .ZN(n24376) );
  INV_X1 U28847 ( .A(n24376), .ZN(p_wishbone_bd_ram_n25904) );
  INV_X1 U28848 ( .A(n64040), .ZN(n24378) );
  INV_X1 U28849 ( .A(n24378), .ZN(p_wishbone_bd_ram_n25903) );
  INV_X1 U28850 ( .A(n64039), .ZN(n24380) );
  INV_X1 U28851 ( .A(n24380), .ZN(p_wishbone_bd_ram_n25902) );
  INV_X1 U28852 ( .A(n64038), .ZN(n24382) );
  INV_X1 U28853 ( .A(n24382), .ZN(p_wishbone_bd_ram_n25901) );
  INV_X1 U28854 ( .A(n64037), .ZN(n24384) );
  INV_X1 U28855 ( .A(n24384), .ZN(p_wishbone_bd_ram_n25900) );
  INV_X1 U28856 ( .A(n64036), .ZN(n24386) );
  INV_X1 U28857 ( .A(n24386), .ZN(p_wishbone_bd_ram_n25899) );
  INV_X1 U28858 ( .A(n64035), .ZN(n24388) );
  INV_X1 U28859 ( .A(n24388), .ZN(p_wishbone_bd_ram_n25898) );
  INV_X1 U28860 ( .A(n64034), .ZN(n24390) );
  INV_X1 U28861 ( .A(n24390), .ZN(p_wishbone_bd_ram_n25897) );
  INV_X1 U28862 ( .A(n64033), .ZN(n24392) );
  INV_X1 U28863 ( .A(n24392), .ZN(p_wishbone_bd_ram_n25896) );
  INV_X1 U28864 ( .A(n64032), .ZN(n24394) );
  INV_X1 U28865 ( .A(n24394), .ZN(p_wishbone_bd_ram_n25895) );
  INV_X1 U28866 ( .A(n64031), .ZN(n24396) );
  INV_X1 U28867 ( .A(n24396), .ZN(p_wishbone_bd_ram_n25894) );
  INV_X1 U28868 ( .A(n64030), .ZN(n24398) );
  INV_X1 U28869 ( .A(n24398), .ZN(p_wishbone_bd_ram_n25893) );
  INV_X1 U28870 ( .A(n64029), .ZN(n24400) );
  INV_X1 U28871 ( .A(n24400), .ZN(p_wishbone_bd_ram_n25892) );
  INV_X1 U28872 ( .A(n64028), .ZN(n24402) );
  INV_X1 U28873 ( .A(n24402), .ZN(p_wishbone_bd_ram_n25891) );
  INV_X1 U28874 ( .A(n64027), .ZN(n24404) );
  INV_X1 U28875 ( .A(n24404), .ZN(p_wishbone_bd_ram_n25890) );
  INV_X1 U28876 ( .A(n64026), .ZN(n24406) );
  INV_X1 U28877 ( .A(n24406), .ZN(p_wishbone_bd_ram_n25889) );
  INV_X1 U28878 ( .A(n64025), .ZN(n24408) );
  INV_X1 U28879 ( .A(n24408), .ZN(p_wishbone_bd_ram_n25888) );
  INV_X1 U28880 ( .A(n64024), .ZN(n24410) );
  INV_X1 U28881 ( .A(n24410), .ZN(p_wishbone_bd_ram_n25887) );
  INV_X1 U28882 ( .A(n64023), .ZN(n24412) );
  INV_X1 U28883 ( .A(n24412), .ZN(p_wishbone_bd_ram_n25886) );
  INV_X1 U28884 ( .A(n64022), .ZN(n24414) );
  INV_X1 U28885 ( .A(n24414), .ZN(p_wishbone_bd_ram_n25885) );
  INV_X1 U28886 ( .A(n64021), .ZN(n24416) );
  INV_X1 U28887 ( .A(n24416), .ZN(p_wishbone_bd_ram_n25884) );
  INV_X1 U28888 ( .A(n64020), .ZN(n24418) );
  INV_X1 U28889 ( .A(n24418), .ZN(p_wishbone_bd_ram_n25883) );
  INV_X1 U28890 ( .A(n64019), .ZN(n24420) );
  INV_X1 U28891 ( .A(n24420), .ZN(p_wishbone_bd_ram_n25882) );
  INV_X1 U28892 ( .A(n64018), .ZN(n24422) );
  INV_X1 U28893 ( .A(n24422), .ZN(p_wishbone_bd_ram_n25881) );
  INV_X1 U28894 ( .A(n64017), .ZN(n24424) );
  INV_X1 U28895 ( .A(n24424), .ZN(p_wishbone_bd_ram_n25880) );
  INV_X1 U28896 ( .A(n64016), .ZN(n24426) );
  INV_X1 U28897 ( .A(n24426), .ZN(p_wishbone_bd_ram_n25879) );
  INV_X1 U28898 ( .A(n64015), .ZN(n24428) );
  INV_X1 U28899 ( .A(n24428), .ZN(p_wishbone_bd_ram_n25878) );
  INV_X1 U28900 ( .A(n64014), .ZN(n24430) );
  INV_X1 U28901 ( .A(n24430), .ZN(p_wishbone_bd_ram_n25877) );
  INV_X1 U28902 ( .A(n64013), .ZN(n24432) );
  INV_X1 U28903 ( .A(n24432), .ZN(p_wishbone_bd_ram_n25876) );
  INV_X1 U28904 ( .A(n64012), .ZN(n24434) );
  INV_X1 U28905 ( .A(n24434), .ZN(p_wishbone_bd_ram_n25875) );
  INV_X1 U28906 ( .A(n64011), .ZN(n24436) );
  INV_X1 U28907 ( .A(n24436), .ZN(p_wishbone_bd_ram_n25874) );
  INV_X1 U28908 ( .A(n64010), .ZN(n24438) );
  INV_X1 U28909 ( .A(n24438), .ZN(p_wishbone_bd_ram_n25873) );
  INV_X1 U28910 ( .A(n64009), .ZN(n24440) );
  INV_X1 U28911 ( .A(n24440), .ZN(p_wishbone_bd_ram_n25872) );
  INV_X1 U28912 ( .A(n64008), .ZN(n24442) );
  INV_X1 U28913 ( .A(n24442), .ZN(p_wishbone_bd_ram_n25871) );
  INV_X1 U28914 ( .A(n64007), .ZN(n24444) );
  INV_X1 U28915 ( .A(n24444), .ZN(p_wishbone_bd_ram_n25870) );
  INV_X1 U28916 ( .A(n64006), .ZN(n24446) );
  INV_X1 U28917 ( .A(n24446), .ZN(p_wishbone_bd_ram_n25869) );
  INV_X1 U28918 ( .A(n64005), .ZN(n24448) );
  INV_X1 U28919 ( .A(n24448), .ZN(p_wishbone_bd_ram_n25868) );
  INV_X1 U28920 ( .A(n64004), .ZN(n24450) );
  INV_X1 U28921 ( .A(n24450), .ZN(p_wishbone_bd_ram_n25867) );
  INV_X1 U28922 ( .A(n64003), .ZN(n24452) );
  INV_X1 U28923 ( .A(n24452), .ZN(p_wishbone_bd_ram_n25866) );
  INV_X1 U28924 ( .A(n64002), .ZN(n24454) );
  INV_X1 U28925 ( .A(n24454), .ZN(p_wishbone_bd_ram_n25865) );
  INV_X1 U28926 ( .A(n64001), .ZN(n24456) );
  INV_X1 U28927 ( .A(n24456), .ZN(p_wishbone_bd_ram_n25864) );
  INV_X1 U28928 ( .A(n64000), .ZN(n24458) );
  INV_X1 U28929 ( .A(n24458), .ZN(p_wishbone_bd_ram_n25863) );
  INV_X1 U28930 ( .A(n63999), .ZN(n24460) );
  INV_X1 U28931 ( .A(n24460), .ZN(p_wishbone_bd_ram_n25862) );
  INV_X1 U28932 ( .A(n63998), .ZN(n24462) );
  INV_X1 U28933 ( .A(n24462), .ZN(p_wishbone_bd_ram_n25861) );
  INV_X1 U28934 ( .A(n63997), .ZN(n24464) );
  INV_X1 U28935 ( .A(n24464), .ZN(p_wishbone_bd_ram_n25860) );
  INV_X1 U28936 ( .A(n63996), .ZN(n24466) );
  INV_X1 U28937 ( .A(n24466), .ZN(p_wishbone_bd_ram_n25859) );
  INV_X1 U28938 ( .A(n63995), .ZN(n24468) );
  INV_X1 U28939 ( .A(n24468), .ZN(p_wishbone_bd_ram_n25858) );
  INV_X1 U28940 ( .A(n63994), .ZN(n24470) );
  INV_X1 U28941 ( .A(n24470), .ZN(p_wishbone_bd_ram_n25857) );
  INV_X1 U28942 ( .A(n63993), .ZN(n24472) );
  INV_X1 U28943 ( .A(n24472), .ZN(p_wishbone_bd_ram_n25856) );
  INV_X1 U28944 ( .A(n63992), .ZN(n24474) );
  INV_X1 U28945 ( .A(n24474), .ZN(p_wishbone_bd_ram_n25855) );
  INV_X1 U28946 ( .A(n63991), .ZN(n24476) );
  INV_X1 U28947 ( .A(n24476), .ZN(p_wishbone_bd_ram_n25854) );
  INV_X1 U28948 ( .A(n63990), .ZN(n24478) );
  INV_X1 U28949 ( .A(n24478), .ZN(p_wishbone_bd_ram_n25853) );
  INV_X1 U28950 ( .A(n63989), .ZN(n24480) );
  INV_X1 U28951 ( .A(n24480), .ZN(p_wishbone_bd_ram_n25852) );
  INV_X1 U28952 ( .A(n63988), .ZN(n24482) );
  INV_X1 U28953 ( .A(n24482), .ZN(p_wishbone_bd_ram_n25851) );
  INV_X1 U28954 ( .A(n63987), .ZN(n24484) );
  INV_X1 U28955 ( .A(n24484), .ZN(p_wishbone_bd_ram_n25850) );
  INV_X1 U28956 ( .A(n63986), .ZN(n24486) );
  INV_X1 U28957 ( .A(n24486), .ZN(p_wishbone_bd_ram_n25849) );
  INV_X1 U28958 ( .A(n63985), .ZN(n24488) );
  INV_X1 U28959 ( .A(n24488), .ZN(p_wishbone_bd_ram_n25848) );
  INV_X1 U28960 ( .A(n63984), .ZN(n24490) );
  INV_X1 U28961 ( .A(n24490), .ZN(p_wishbone_bd_ram_n25847) );
  INV_X1 U28962 ( .A(n63983), .ZN(n24492) );
  INV_X1 U28963 ( .A(n24492), .ZN(p_wishbone_bd_ram_n25846) );
  INV_X1 U28964 ( .A(n63982), .ZN(n24494) );
  INV_X1 U28965 ( .A(n24494), .ZN(p_wishbone_bd_ram_n25845) );
  INV_X1 U28966 ( .A(n63981), .ZN(n24496) );
  INV_X1 U28967 ( .A(n24496), .ZN(p_wishbone_bd_ram_n25844) );
  INV_X1 U28968 ( .A(n63980), .ZN(n24498) );
  INV_X1 U28969 ( .A(n24498), .ZN(p_wishbone_bd_ram_n25843) );
  INV_X1 U28970 ( .A(n63979), .ZN(n24500) );
  INV_X1 U28971 ( .A(n24500), .ZN(p_wishbone_bd_ram_n25842) );
  INV_X1 U28972 ( .A(n63978), .ZN(n24502) );
  INV_X1 U28973 ( .A(n24502), .ZN(p_wishbone_bd_ram_n25841) );
  INV_X1 U28974 ( .A(n63977), .ZN(n24504) );
  INV_X1 U28975 ( .A(n24504), .ZN(p_wishbone_bd_ram_n25840) );
  INV_X1 U28976 ( .A(n63976), .ZN(n24506) );
  INV_X1 U28977 ( .A(n24506), .ZN(p_wishbone_bd_ram_n25839) );
  INV_X1 U28978 ( .A(n63975), .ZN(n24508) );
  INV_X1 U28979 ( .A(n24508), .ZN(p_wishbone_bd_ram_n25838) );
  INV_X1 U28980 ( .A(n63974), .ZN(n24510) );
  INV_X1 U28981 ( .A(n24510), .ZN(p_wishbone_bd_ram_n25837) );
  INV_X1 U28982 ( .A(n63973), .ZN(n24512) );
  INV_X1 U28983 ( .A(n24512), .ZN(p_wishbone_bd_ram_n25836) );
  INV_X1 U28984 ( .A(n63972), .ZN(n24514) );
  INV_X1 U28985 ( .A(n24514), .ZN(p_wishbone_bd_ram_n25835) );
  INV_X1 U28986 ( .A(n63971), .ZN(n24516) );
  INV_X1 U28987 ( .A(n24516), .ZN(p_wishbone_bd_ram_n25834) );
  INV_X1 U28988 ( .A(n63970), .ZN(n24518) );
  INV_X1 U28989 ( .A(n24518), .ZN(p_wishbone_bd_ram_n25833) );
  INV_X1 U28990 ( .A(n63969), .ZN(n24520) );
  INV_X1 U28991 ( .A(n24520), .ZN(p_wishbone_bd_ram_n25832) );
  INV_X1 U28992 ( .A(n63968), .ZN(n24522) );
  INV_X1 U28993 ( .A(n24522), .ZN(p_wishbone_bd_ram_n25831) );
  INV_X1 U28994 ( .A(n63967), .ZN(n24524) );
  INV_X1 U28995 ( .A(n24524), .ZN(p_wishbone_bd_ram_n25830) );
  INV_X1 U28996 ( .A(n63966), .ZN(n24526) );
  INV_X1 U28997 ( .A(n24526), .ZN(p_wishbone_bd_ram_n25829) );
  INV_X1 U28998 ( .A(n63965), .ZN(n24528) );
  INV_X1 U28999 ( .A(n24528), .ZN(p_wishbone_bd_ram_n25828) );
  INV_X1 U29000 ( .A(n63964), .ZN(n24530) );
  INV_X1 U29001 ( .A(n24530), .ZN(p_wishbone_bd_ram_n25827) );
  INV_X1 U29002 ( .A(n63963), .ZN(n24532) );
  INV_X1 U29003 ( .A(n24532), .ZN(p_wishbone_bd_ram_n25826) );
  INV_X1 U29004 ( .A(n63962), .ZN(n24534) );
  INV_X1 U29005 ( .A(n24534), .ZN(p_wishbone_bd_ram_n25825) );
  INV_X1 U29006 ( .A(n63961), .ZN(n24536) );
  INV_X1 U29007 ( .A(n24536), .ZN(p_wishbone_bd_ram_n25824) );
  INV_X1 U29008 ( .A(n63960), .ZN(n24538) );
  INV_X1 U29009 ( .A(n24538), .ZN(p_wishbone_bd_ram_n25823) );
  INV_X1 U29010 ( .A(n63959), .ZN(n24540) );
  INV_X1 U29011 ( .A(n24540), .ZN(p_wishbone_bd_ram_n25822) );
  INV_X1 U29012 ( .A(n63958), .ZN(n24542) );
  INV_X1 U29013 ( .A(n24542), .ZN(p_wishbone_bd_ram_n25821) );
  INV_X1 U29014 ( .A(n63957), .ZN(n24544) );
  INV_X1 U29015 ( .A(n24544), .ZN(p_wishbone_bd_ram_n25820) );
  INV_X1 U29016 ( .A(n63956), .ZN(n24546) );
  INV_X1 U29017 ( .A(n24546), .ZN(p_wishbone_bd_ram_n25819) );
  INV_X1 U29018 ( .A(n63955), .ZN(n24548) );
  INV_X1 U29019 ( .A(n24548), .ZN(p_wishbone_bd_ram_n25818) );
  INV_X1 U29020 ( .A(n63954), .ZN(n24550) );
  INV_X1 U29021 ( .A(n24550), .ZN(p_wishbone_bd_ram_n25817) );
  INV_X1 U29022 ( .A(n63953), .ZN(n24552) );
  INV_X1 U29023 ( .A(n24552), .ZN(p_wishbone_bd_ram_n25816) );
  INV_X1 U29024 ( .A(n63952), .ZN(n24554) );
  INV_X1 U29025 ( .A(n24554), .ZN(p_wishbone_bd_ram_n25815) );
  INV_X1 U29026 ( .A(n63951), .ZN(n24556) );
  INV_X1 U29027 ( .A(n24556), .ZN(p_wishbone_bd_ram_n25814) );
  INV_X1 U29028 ( .A(n63950), .ZN(n24558) );
  INV_X1 U29029 ( .A(n24558), .ZN(p_wishbone_bd_ram_n25813) );
  INV_X1 U29030 ( .A(n63949), .ZN(n24560) );
  INV_X1 U29031 ( .A(n24560), .ZN(p_wishbone_bd_ram_n25812) );
  INV_X1 U29032 ( .A(n63948), .ZN(n24562) );
  INV_X1 U29033 ( .A(n24562), .ZN(p_wishbone_bd_ram_n25811) );
  INV_X1 U29034 ( .A(n63947), .ZN(n24564) );
  INV_X1 U29035 ( .A(n24564), .ZN(p_wishbone_bd_ram_n25810) );
  INV_X1 U29036 ( .A(n63946), .ZN(n24566) );
  INV_X1 U29037 ( .A(n24566), .ZN(p_wishbone_bd_ram_n25809) );
  INV_X1 U29038 ( .A(n63945), .ZN(n24568) );
  INV_X1 U29039 ( .A(n24568), .ZN(p_wishbone_bd_ram_n25808) );
  INV_X1 U29040 ( .A(n63944), .ZN(n24570) );
  INV_X1 U29041 ( .A(n24570), .ZN(p_wishbone_bd_ram_n25807) );
  INV_X1 U29042 ( .A(n63943), .ZN(n24572) );
  INV_X1 U29043 ( .A(n24572), .ZN(p_wishbone_bd_ram_n25806) );
  INV_X1 U29044 ( .A(n63942), .ZN(n24574) );
  INV_X1 U29045 ( .A(n24574), .ZN(p_wishbone_bd_ram_n25805) );
  INV_X1 U29046 ( .A(n63941), .ZN(n24576) );
  INV_X1 U29047 ( .A(n24576), .ZN(p_wishbone_bd_ram_n25804) );
  INV_X1 U29048 ( .A(n63940), .ZN(n24578) );
  INV_X1 U29049 ( .A(n24578), .ZN(p_wishbone_bd_ram_n25803) );
  INV_X1 U29050 ( .A(n63939), .ZN(n24580) );
  INV_X1 U29051 ( .A(n24580), .ZN(p_wishbone_bd_ram_n25802) );
  INV_X1 U29052 ( .A(n63938), .ZN(n24582) );
  INV_X1 U29053 ( .A(n24582), .ZN(p_wishbone_bd_ram_n25801) );
  INV_X1 U29054 ( .A(n63937), .ZN(n24584) );
  INV_X1 U29055 ( .A(n24584), .ZN(p_wishbone_bd_ram_n25800) );
  INV_X1 U29056 ( .A(n63936), .ZN(n24586) );
  INV_X1 U29057 ( .A(n24586), .ZN(p_wishbone_bd_ram_n25799) );
  INV_X1 U29058 ( .A(n63935), .ZN(n24588) );
  INV_X1 U29059 ( .A(n24588), .ZN(p_wishbone_bd_ram_n25798) );
  INV_X1 U29060 ( .A(n63934), .ZN(n24590) );
  INV_X1 U29061 ( .A(n24590), .ZN(p_wishbone_bd_ram_n25797) );
  INV_X1 U29062 ( .A(n63933), .ZN(n24592) );
  INV_X1 U29063 ( .A(n24592), .ZN(p_wishbone_bd_ram_n25796) );
  INV_X1 U29064 ( .A(n63932), .ZN(n24594) );
  INV_X1 U29065 ( .A(n24594), .ZN(p_wishbone_bd_ram_n25795) );
  INV_X1 U29066 ( .A(n63931), .ZN(n24596) );
  INV_X1 U29067 ( .A(n24596), .ZN(p_wishbone_bd_ram_n25794) );
  INV_X1 U29068 ( .A(n63930), .ZN(n24598) );
  INV_X1 U29069 ( .A(n24598), .ZN(p_wishbone_bd_ram_n25793) );
  INV_X1 U29070 ( .A(n63929), .ZN(n24600) );
  INV_X1 U29071 ( .A(n24600), .ZN(p_wishbone_bd_ram_n25792) );
  INV_X1 U29072 ( .A(n63928), .ZN(n24602) );
  INV_X1 U29073 ( .A(n24602), .ZN(p_wishbone_bd_ram_n25791) );
  INV_X1 U29074 ( .A(n63927), .ZN(n24604) );
  INV_X1 U29075 ( .A(n24604), .ZN(p_wishbone_bd_ram_n25790) );
  INV_X1 U29076 ( .A(n63926), .ZN(n24606) );
  INV_X1 U29077 ( .A(n24606), .ZN(p_wishbone_bd_ram_n25789) );
  INV_X1 U29078 ( .A(n63925), .ZN(n24608) );
  INV_X1 U29079 ( .A(n24608), .ZN(p_wishbone_bd_ram_n25788) );
  INV_X1 U29080 ( .A(n63924), .ZN(n24610) );
  INV_X1 U29081 ( .A(n24610), .ZN(p_wishbone_bd_ram_n25787) );
  INV_X1 U29082 ( .A(n63923), .ZN(n24612) );
  INV_X1 U29083 ( .A(n24612), .ZN(p_wishbone_bd_ram_n25786) );
  INV_X1 U29084 ( .A(n63922), .ZN(n24614) );
  INV_X1 U29085 ( .A(n24614), .ZN(p_wishbone_bd_ram_n25785) );
  INV_X1 U29086 ( .A(n63921), .ZN(n24616) );
  INV_X1 U29087 ( .A(n24616), .ZN(p_wishbone_bd_ram_n25784) );
  INV_X1 U29088 ( .A(n63920), .ZN(n24618) );
  INV_X1 U29089 ( .A(n24618), .ZN(p_wishbone_bd_ram_n25783) );
  INV_X1 U29090 ( .A(n63919), .ZN(n24620) );
  INV_X1 U29091 ( .A(n24620), .ZN(p_wishbone_bd_ram_n25782) );
  INV_X1 U29092 ( .A(n63918), .ZN(n24622) );
  INV_X1 U29093 ( .A(n24622), .ZN(p_wishbone_bd_ram_n25781) );
  INV_X1 U29094 ( .A(n63917), .ZN(n24624) );
  INV_X1 U29095 ( .A(n24624), .ZN(p_wishbone_bd_ram_n25780) );
  INV_X1 U29096 ( .A(n63916), .ZN(n24626) );
  INV_X1 U29097 ( .A(n24626), .ZN(p_wishbone_bd_ram_n25779) );
  INV_X1 U29098 ( .A(n63915), .ZN(n24628) );
  INV_X1 U29099 ( .A(n24628), .ZN(p_wishbone_bd_ram_n25778) );
  INV_X1 U29100 ( .A(n63914), .ZN(n24630) );
  INV_X1 U29101 ( .A(n24630), .ZN(p_wishbone_bd_ram_n25777) );
  INV_X1 U29102 ( .A(n63913), .ZN(n24632) );
  INV_X1 U29103 ( .A(n24632), .ZN(p_wishbone_bd_ram_n25776) );
  INV_X1 U29104 ( .A(n63912), .ZN(n24634) );
  INV_X1 U29105 ( .A(n24634), .ZN(p_wishbone_bd_ram_n25775) );
  INV_X1 U29106 ( .A(n63911), .ZN(n24636) );
  INV_X1 U29107 ( .A(n24636), .ZN(p_wishbone_bd_ram_n25774) );
  INV_X1 U29108 ( .A(n63910), .ZN(n24638) );
  INV_X1 U29109 ( .A(n24638), .ZN(p_wishbone_bd_ram_n25773) );
  INV_X1 U29110 ( .A(n63909), .ZN(n24640) );
  INV_X1 U29111 ( .A(n24640), .ZN(p_wishbone_bd_ram_n25772) );
  INV_X1 U29112 ( .A(n63908), .ZN(n24642) );
  INV_X1 U29113 ( .A(n24642), .ZN(p_wishbone_bd_ram_n25771) );
  INV_X1 U29114 ( .A(n63907), .ZN(n24644) );
  INV_X1 U29115 ( .A(n24644), .ZN(p_wishbone_bd_ram_n25770) );
  INV_X1 U29116 ( .A(n63906), .ZN(n24646) );
  INV_X1 U29117 ( .A(n24646), .ZN(p_wishbone_bd_ram_n25769) );
  INV_X1 U29118 ( .A(n63905), .ZN(n24648) );
  INV_X1 U29119 ( .A(n24648), .ZN(p_wishbone_bd_ram_n25768) );
  INV_X1 U29120 ( .A(n63904), .ZN(n24650) );
  INV_X1 U29121 ( .A(n24650), .ZN(p_wishbone_bd_ram_n25767) );
  INV_X1 U29122 ( .A(n63903), .ZN(n24652) );
  INV_X1 U29123 ( .A(n24652), .ZN(p_wishbone_bd_ram_n25766) );
  INV_X1 U29124 ( .A(n63902), .ZN(n24654) );
  INV_X1 U29125 ( .A(n24654), .ZN(p_wishbone_bd_ram_n25765) );
  INV_X1 U29126 ( .A(n63901), .ZN(n24656) );
  INV_X1 U29127 ( .A(n24656), .ZN(p_wishbone_bd_ram_n25764) );
  INV_X1 U29128 ( .A(n63900), .ZN(n24658) );
  INV_X1 U29129 ( .A(n24658), .ZN(p_wishbone_bd_ram_n25763) );
  INV_X1 U29130 ( .A(n63899), .ZN(n24660) );
  INV_X1 U29131 ( .A(n24660), .ZN(p_wishbone_bd_ram_n25762) );
  INV_X1 U29132 ( .A(n63898), .ZN(n24662) );
  INV_X1 U29133 ( .A(n24662), .ZN(p_wishbone_bd_ram_n25761) );
  INV_X1 U29134 ( .A(n63897), .ZN(n24664) );
  INV_X1 U29135 ( .A(n24664), .ZN(p_wishbone_bd_ram_n25760) );
  INV_X1 U29136 ( .A(n63896), .ZN(n24666) );
  INV_X1 U29137 ( .A(n24666), .ZN(p_wishbone_bd_ram_n25759) );
  INV_X1 U29138 ( .A(n63895), .ZN(n24668) );
  INV_X1 U29139 ( .A(n24668), .ZN(p_wishbone_bd_ram_n25758) );
  INV_X1 U29140 ( .A(n63894), .ZN(n24670) );
  INV_X1 U29141 ( .A(n24670), .ZN(p_wishbone_bd_ram_n25757) );
  INV_X1 U29142 ( .A(n63893), .ZN(n24672) );
  INV_X1 U29143 ( .A(n24672), .ZN(p_wishbone_bd_ram_n25756) );
  INV_X1 U29144 ( .A(n63892), .ZN(n24674) );
  INV_X1 U29145 ( .A(n24674), .ZN(p_wishbone_bd_ram_n25755) );
  INV_X1 U29146 ( .A(n63891), .ZN(n24676) );
  INV_X1 U29147 ( .A(n24676), .ZN(p_wishbone_bd_ram_n25754) );
  INV_X1 U29148 ( .A(n63890), .ZN(n24678) );
  INV_X1 U29149 ( .A(n24678), .ZN(p_wishbone_bd_ram_n25753) );
  INV_X1 U29150 ( .A(n63889), .ZN(n24680) );
  INV_X1 U29151 ( .A(n24680), .ZN(p_wishbone_bd_ram_n25752) );
  INV_X1 U29152 ( .A(n63888), .ZN(n24682) );
  INV_X1 U29153 ( .A(n24682), .ZN(p_wishbone_bd_ram_n25751) );
  INV_X1 U29154 ( .A(n63887), .ZN(n24684) );
  INV_X1 U29155 ( .A(n24684), .ZN(p_wishbone_bd_ram_n25750) );
  INV_X1 U29156 ( .A(n63886), .ZN(n24686) );
  INV_X1 U29157 ( .A(n24686), .ZN(p_wishbone_bd_ram_n25749) );
  INV_X1 U29158 ( .A(n63885), .ZN(n24688) );
  INV_X1 U29159 ( .A(n24688), .ZN(p_wishbone_bd_ram_n25748) );
  INV_X1 U29160 ( .A(n63884), .ZN(n24690) );
  INV_X1 U29161 ( .A(n24690), .ZN(p_wishbone_bd_ram_n25747) );
  INV_X1 U29162 ( .A(n63883), .ZN(n24692) );
  INV_X1 U29163 ( .A(n24692), .ZN(p_wishbone_bd_ram_n25746) );
  INV_X1 U29164 ( .A(n63882), .ZN(n24694) );
  INV_X1 U29165 ( .A(n24694), .ZN(p_wishbone_bd_ram_n25745) );
  INV_X1 U29166 ( .A(n63881), .ZN(n24696) );
  INV_X1 U29167 ( .A(n24696), .ZN(p_wishbone_bd_ram_n25744) );
  INV_X1 U29168 ( .A(n63880), .ZN(n24698) );
  INV_X1 U29169 ( .A(n24698), .ZN(p_wishbone_bd_ram_n25743) );
  INV_X1 U29170 ( .A(n63879), .ZN(n24700) );
  INV_X1 U29171 ( .A(n24700), .ZN(p_wishbone_bd_ram_n25742) );
  INV_X1 U29172 ( .A(n63878), .ZN(n24702) );
  INV_X1 U29173 ( .A(n24702), .ZN(p_wishbone_bd_ram_n25741) );
  INV_X1 U29174 ( .A(n63877), .ZN(n24704) );
  INV_X1 U29175 ( .A(n24704), .ZN(p_wishbone_bd_ram_n25740) );
  INV_X1 U29176 ( .A(n63876), .ZN(n24706) );
  INV_X1 U29177 ( .A(n24706), .ZN(p_wishbone_bd_ram_n25739) );
  INV_X1 U29178 ( .A(n63875), .ZN(n24708) );
  INV_X1 U29179 ( .A(n24708), .ZN(p_wishbone_bd_ram_n25738) );
  INV_X1 U29180 ( .A(n63874), .ZN(n24710) );
  INV_X1 U29181 ( .A(n24710), .ZN(p_wishbone_bd_ram_n25737) );
  INV_X1 U29182 ( .A(n63873), .ZN(n24712) );
  INV_X1 U29183 ( .A(n24712), .ZN(p_wishbone_bd_ram_n25736) );
  INV_X1 U29184 ( .A(n63872), .ZN(n24714) );
  INV_X1 U29185 ( .A(n24714), .ZN(p_wishbone_bd_ram_n25735) );
  INV_X1 U29186 ( .A(n63871), .ZN(n24716) );
  INV_X1 U29187 ( .A(n24716), .ZN(p_wishbone_bd_ram_n25734) );
  INV_X1 U29188 ( .A(n63870), .ZN(n24718) );
  INV_X1 U29189 ( .A(n24718), .ZN(p_wishbone_bd_ram_n25733) );
  INV_X1 U29190 ( .A(n63869), .ZN(n24720) );
  INV_X1 U29191 ( .A(n24720), .ZN(p_wishbone_bd_ram_n25732) );
  INV_X1 U29192 ( .A(n63868), .ZN(n24722) );
  INV_X1 U29193 ( .A(n24722), .ZN(p_wishbone_bd_ram_n25731) );
  INV_X1 U29194 ( .A(n63867), .ZN(n24724) );
  INV_X1 U29195 ( .A(n24724), .ZN(p_wishbone_bd_ram_n25730) );
  INV_X1 U29196 ( .A(n63866), .ZN(n24726) );
  INV_X1 U29197 ( .A(n24726), .ZN(p_wishbone_bd_ram_n25729) );
  INV_X1 U29198 ( .A(n63865), .ZN(n24728) );
  INV_X1 U29199 ( .A(n24728), .ZN(p_wishbone_bd_ram_n25728) );
  INV_X1 U29200 ( .A(n63864), .ZN(n24730) );
  INV_X1 U29201 ( .A(n24730), .ZN(p_wishbone_bd_ram_n25727) );
  INV_X1 U29202 ( .A(n63863), .ZN(n24732) );
  INV_X1 U29203 ( .A(n24732), .ZN(p_wishbone_bd_ram_n25726) );
  INV_X1 U29204 ( .A(n63862), .ZN(n24734) );
  INV_X1 U29205 ( .A(n24734), .ZN(p_wishbone_bd_ram_n25725) );
  INV_X1 U29206 ( .A(n63861), .ZN(n24736) );
  INV_X1 U29207 ( .A(n24736), .ZN(p_wishbone_bd_ram_n25724) );
  INV_X1 U29208 ( .A(n63860), .ZN(n24738) );
  INV_X1 U29209 ( .A(n24738), .ZN(p_wishbone_bd_ram_n25723) );
  INV_X1 U29210 ( .A(n63859), .ZN(n24740) );
  INV_X1 U29211 ( .A(n24740), .ZN(p_wishbone_bd_ram_n25722) );
  INV_X1 U29212 ( .A(n63858), .ZN(n24742) );
  INV_X1 U29213 ( .A(n24742), .ZN(p_wishbone_bd_ram_n25721) );
  INV_X1 U29214 ( .A(n63857), .ZN(n24744) );
  INV_X1 U29215 ( .A(n24744), .ZN(p_wishbone_bd_ram_n25720) );
  INV_X1 U29216 ( .A(n63856), .ZN(n24746) );
  INV_X1 U29217 ( .A(n24746), .ZN(p_wishbone_bd_ram_n25719) );
  INV_X1 U29218 ( .A(n63855), .ZN(n24748) );
  INV_X1 U29219 ( .A(n24748), .ZN(p_wishbone_bd_ram_n25718) );
  INV_X1 U29220 ( .A(n63854), .ZN(n24750) );
  INV_X1 U29221 ( .A(n24750), .ZN(p_wishbone_bd_ram_n25717) );
  INV_X1 U29222 ( .A(n63853), .ZN(n24752) );
  INV_X1 U29223 ( .A(n24752), .ZN(p_wishbone_bd_ram_n25716) );
  INV_X1 U29224 ( .A(n63852), .ZN(n24754) );
  INV_X1 U29225 ( .A(n24754), .ZN(p_wishbone_bd_ram_n25715) );
  INV_X1 U29226 ( .A(n63851), .ZN(n24756) );
  INV_X1 U29227 ( .A(n24756), .ZN(p_wishbone_bd_ram_n25714) );
  INV_X1 U29228 ( .A(n63850), .ZN(n24758) );
  INV_X1 U29229 ( .A(n24758), .ZN(p_wishbone_bd_ram_n25713) );
  INV_X1 U29230 ( .A(n63849), .ZN(n24760) );
  INV_X1 U29231 ( .A(n24760), .ZN(p_wishbone_bd_ram_n25712) );
  INV_X1 U29232 ( .A(n63848), .ZN(n24762) );
  INV_X1 U29233 ( .A(n24762), .ZN(p_wishbone_bd_ram_n25711) );
  INV_X1 U29234 ( .A(n63847), .ZN(n24764) );
  INV_X1 U29235 ( .A(n24764), .ZN(p_wishbone_bd_ram_n25710) );
  INV_X1 U29236 ( .A(n63846), .ZN(n24766) );
  INV_X1 U29237 ( .A(n24766), .ZN(p_wishbone_bd_ram_n25709) );
  INV_X1 U29238 ( .A(n63845), .ZN(n24768) );
  INV_X1 U29239 ( .A(n24768), .ZN(p_wishbone_bd_ram_n25708) );
  INV_X1 U29240 ( .A(n63844), .ZN(n24770) );
  INV_X1 U29241 ( .A(n24770), .ZN(p_wishbone_bd_ram_n25707) );
  INV_X1 U29242 ( .A(n63843), .ZN(n24772) );
  INV_X1 U29243 ( .A(n24772), .ZN(p_wishbone_bd_ram_n25706) );
  INV_X1 U29244 ( .A(n63842), .ZN(n24774) );
  INV_X1 U29245 ( .A(n24774), .ZN(p_wishbone_bd_ram_n25705) );
  INV_X1 U29246 ( .A(n63841), .ZN(n24776) );
  INV_X1 U29247 ( .A(n24776), .ZN(p_wishbone_bd_ram_n25704) );
  INV_X1 U29248 ( .A(n63840), .ZN(n24778) );
  INV_X1 U29249 ( .A(n24778), .ZN(p_wishbone_bd_ram_n25703) );
  INV_X1 U29250 ( .A(n63839), .ZN(n24780) );
  INV_X1 U29251 ( .A(n24780), .ZN(p_wishbone_bd_ram_n25702) );
  INV_X1 U29252 ( .A(n63838), .ZN(n24782) );
  INV_X1 U29253 ( .A(n24782), .ZN(p_wishbone_bd_ram_n25701) );
  INV_X1 U29254 ( .A(n63837), .ZN(n24784) );
  INV_X1 U29255 ( .A(n24784), .ZN(p_wishbone_bd_ram_n25700) );
  INV_X1 U29256 ( .A(n63836), .ZN(n24786) );
  INV_X1 U29257 ( .A(n24786), .ZN(p_wishbone_bd_ram_n25699) );
  INV_X1 U29258 ( .A(n63835), .ZN(n24788) );
  INV_X1 U29259 ( .A(n24788), .ZN(p_wishbone_bd_ram_n25698) );
  INV_X1 U29260 ( .A(n63834), .ZN(n24790) );
  INV_X1 U29261 ( .A(n24790), .ZN(p_wishbone_bd_ram_n25697) );
  INV_X1 U29262 ( .A(n63833), .ZN(n24792) );
  INV_X1 U29263 ( .A(n24792), .ZN(p_wishbone_bd_ram_n25696) );
  INV_X1 U29264 ( .A(n63832), .ZN(n24794) );
  INV_X1 U29265 ( .A(n24794), .ZN(p_wishbone_bd_ram_n25695) );
  INV_X1 U29266 ( .A(n63831), .ZN(n24796) );
  INV_X1 U29267 ( .A(n24796), .ZN(p_wishbone_bd_ram_n25694) );
  INV_X1 U29268 ( .A(n63830), .ZN(n24798) );
  INV_X1 U29269 ( .A(n24798), .ZN(p_wishbone_bd_ram_n25693) );
  INV_X1 U29270 ( .A(n63829), .ZN(n24800) );
  INV_X1 U29271 ( .A(n24800), .ZN(p_wishbone_bd_ram_n25692) );
  INV_X1 U29272 ( .A(n63828), .ZN(n24802) );
  INV_X1 U29273 ( .A(n24802), .ZN(p_wishbone_bd_ram_n25691) );
  INV_X1 U29274 ( .A(n63827), .ZN(n24804) );
  INV_X1 U29275 ( .A(n24804), .ZN(p_wishbone_bd_ram_n25690) );
  INV_X1 U29276 ( .A(n63826), .ZN(n24806) );
  INV_X1 U29277 ( .A(n24806), .ZN(p_wishbone_bd_ram_n25689) );
  INV_X1 U29278 ( .A(n63825), .ZN(n24808) );
  INV_X1 U29279 ( .A(n24808), .ZN(p_wishbone_bd_ram_n25688) );
  INV_X1 U29280 ( .A(n63824), .ZN(n24810) );
  INV_X1 U29281 ( .A(n24810), .ZN(p_wishbone_bd_ram_n25687) );
  INV_X1 U29282 ( .A(n63823), .ZN(n24812) );
  INV_X1 U29283 ( .A(n24812), .ZN(p_wishbone_bd_ram_n25686) );
  INV_X1 U29284 ( .A(n63822), .ZN(n24814) );
  INV_X1 U29285 ( .A(n24814), .ZN(p_wishbone_bd_ram_n25685) );
  INV_X1 U29286 ( .A(n63821), .ZN(n24816) );
  INV_X1 U29287 ( .A(n24816), .ZN(p_wishbone_bd_ram_n25684) );
  INV_X1 U29288 ( .A(n63820), .ZN(n24818) );
  INV_X1 U29289 ( .A(n24818), .ZN(p_wishbone_bd_ram_n25683) );
  INV_X1 U29290 ( .A(n63819), .ZN(n24820) );
  INV_X1 U29291 ( .A(n24820), .ZN(p_wishbone_bd_ram_n25682) );
  INV_X1 U29292 ( .A(n63818), .ZN(n24822) );
  INV_X1 U29293 ( .A(n24822), .ZN(p_wishbone_bd_ram_n25681) );
  INV_X1 U29294 ( .A(n63817), .ZN(n24824) );
  INV_X1 U29295 ( .A(n24824), .ZN(p_wishbone_bd_ram_n25680) );
  INV_X1 U29296 ( .A(n63816), .ZN(n24826) );
  INV_X1 U29297 ( .A(n24826), .ZN(p_wishbone_bd_ram_n25679) );
  INV_X1 U29298 ( .A(n63815), .ZN(n24828) );
  INV_X1 U29299 ( .A(n24828), .ZN(p_wishbone_bd_ram_n25678) );
  INV_X1 U29300 ( .A(n63814), .ZN(n24830) );
  INV_X1 U29301 ( .A(n24830), .ZN(p_wishbone_bd_ram_n25677) );
  INV_X1 U29302 ( .A(n63813), .ZN(n24832) );
  INV_X1 U29303 ( .A(n24832), .ZN(p_wishbone_bd_ram_n25676) );
  INV_X1 U29304 ( .A(n63812), .ZN(n24834) );
  INV_X1 U29305 ( .A(n24834), .ZN(p_wishbone_bd_ram_n25675) );
  INV_X1 U29306 ( .A(n63811), .ZN(n24836) );
  INV_X1 U29307 ( .A(n24836), .ZN(p_wishbone_bd_ram_n25674) );
  INV_X1 U29308 ( .A(n63810), .ZN(n24838) );
  INV_X1 U29309 ( .A(n24838), .ZN(p_wishbone_bd_ram_n25673) );
  INV_X1 U29310 ( .A(n63809), .ZN(n24840) );
  INV_X1 U29311 ( .A(n24840), .ZN(p_wishbone_bd_ram_n25672) );
  INV_X1 U29312 ( .A(n63808), .ZN(n24842) );
  INV_X1 U29313 ( .A(n24842), .ZN(p_wishbone_bd_ram_n25671) );
  INV_X1 U29314 ( .A(n63807), .ZN(n24844) );
  INV_X1 U29315 ( .A(n24844), .ZN(p_wishbone_bd_ram_n25670) );
  INV_X1 U29316 ( .A(n63806), .ZN(n24846) );
  INV_X1 U29317 ( .A(n24846), .ZN(p_wishbone_bd_ram_n25669) );
  INV_X1 U29318 ( .A(n63805), .ZN(n24848) );
  INV_X1 U29319 ( .A(n24848), .ZN(p_wishbone_bd_ram_n25668) );
  INV_X1 U29320 ( .A(n63804), .ZN(n24850) );
  INV_X1 U29321 ( .A(n24850), .ZN(p_wishbone_bd_ram_n25667) );
  INV_X1 U29322 ( .A(n63803), .ZN(n24852) );
  INV_X1 U29323 ( .A(n24852), .ZN(p_wishbone_bd_ram_n25666) );
  INV_X1 U29324 ( .A(n63802), .ZN(n24854) );
  INV_X1 U29325 ( .A(n24854), .ZN(p_wishbone_bd_ram_n25665) );
  INV_X1 U29326 ( .A(n63801), .ZN(n24856) );
  INV_X1 U29327 ( .A(n24856), .ZN(p_wishbone_bd_ram_n25664) );
  INV_X1 U29328 ( .A(n63800), .ZN(n24858) );
  INV_X1 U29329 ( .A(n24858), .ZN(p_wishbone_bd_ram_n25663) );
  INV_X1 U29330 ( .A(n63799), .ZN(n24860) );
  INV_X1 U29331 ( .A(n24860), .ZN(p_wishbone_bd_ram_n25662) );
  INV_X1 U29332 ( .A(n63798), .ZN(n24862) );
  INV_X1 U29333 ( .A(n24862), .ZN(p_wishbone_bd_ram_n25661) );
  INV_X1 U29334 ( .A(n63797), .ZN(n24864) );
  INV_X1 U29335 ( .A(n24864), .ZN(p_wishbone_bd_ram_n25660) );
  INV_X1 U29336 ( .A(n63796), .ZN(n24866) );
  INV_X1 U29337 ( .A(n24866), .ZN(p_wishbone_bd_ram_n25659) );
  INV_X1 U29338 ( .A(n63795), .ZN(n24868) );
  INV_X1 U29339 ( .A(n24868), .ZN(p_wishbone_bd_ram_n25658) );
  INV_X1 U29340 ( .A(n63794), .ZN(n24870) );
  INV_X1 U29341 ( .A(n24870), .ZN(p_wishbone_bd_ram_n25657) );
  INV_X1 U29342 ( .A(n63793), .ZN(n24872) );
  INV_X1 U29343 ( .A(n24872), .ZN(p_wishbone_bd_ram_n25656) );
  INV_X1 U29344 ( .A(n63792), .ZN(n24874) );
  INV_X1 U29345 ( .A(n24874), .ZN(p_wishbone_bd_ram_n25655) );
  INV_X1 U29346 ( .A(n63791), .ZN(n24876) );
  INV_X1 U29347 ( .A(n24876), .ZN(p_wishbone_bd_ram_n25654) );
  INV_X1 U29348 ( .A(n63790), .ZN(n24878) );
  INV_X1 U29349 ( .A(n24878), .ZN(p_wishbone_bd_ram_n25653) );
  INV_X1 U29350 ( .A(n63789), .ZN(n24880) );
  INV_X1 U29351 ( .A(n24880), .ZN(p_wishbone_bd_ram_n25652) );
  INV_X1 U29352 ( .A(n63788), .ZN(n24882) );
  INV_X1 U29353 ( .A(n24882), .ZN(p_wishbone_bd_ram_n25651) );
  INV_X1 U29354 ( .A(n63787), .ZN(n24884) );
  INV_X1 U29355 ( .A(n24884), .ZN(p_wishbone_bd_ram_n25650) );
  INV_X1 U29356 ( .A(n63786), .ZN(n24886) );
  INV_X1 U29357 ( .A(n24886), .ZN(p_wishbone_bd_ram_n25649) );
  INV_X1 U29358 ( .A(n63785), .ZN(n24888) );
  INV_X1 U29359 ( .A(n24888), .ZN(p_wishbone_bd_ram_n25648) );
  INV_X1 U29360 ( .A(n63784), .ZN(n24890) );
  INV_X1 U29361 ( .A(n24890), .ZN(p_wishbone_bd_ram_n25647) );
  INV_X1 U29362 ( .A(n63783), .ZN(n24892) );
  INV_X1 U29363 ( .A(n24892), .ZN(p_wishbone_bd_ram_n25646) );
  INV_X1 U29364 ( .A(n63782), .ZN(n24894) );
  INV_X1 U29365 ( .A(n24894), .ZN(p_wishbone_bd_ram_n25645) );
  INV_X1 U29366 ( .A(n63781), .ZN(n24896) );
  INV_X1 U29367 ( .A(n24896), .ZN(p_wishbone_bd_ram_n25644) );
  INV_X1 U29368 ( .A(n63780), .ZN(n24898) );
  INV_X1 U29369 ( .A(n24898), .ZN(p_wishbone_bd_ram_n25643) );
  INV_X1 U29370 ( .A(n63779), .ZN(n24900) );
  INV_X1 U29371 ( .A(n24900), .ZN(p_wishbone_bd_ram_n25642) );
  INV_X1 U29372 ( .A(n63778), .ZN(n24902) );
  INV_X1 U29373 ( .A(n24902), .ZN(p_wishbone_bd_ram_n25641) );
  INV_X1 U29374 ( .A(n63777), .ZN(n24904) );
  INV_X1 U29375 ( .A(n24904), .ZN(p_wishbone_bd_ram_n25640) );
  INV_X1 U29376 ( .A(n63776), .ZN(n24906) );
  INV_X1 U29377 ( .A(n24906), .ZN(p_wishbone_bd_ram_n25639) );
  INV_X1 U29378 ( .A(n63775), .ZN(n24908) );
  INV_X1 U29379 ( .A(n24908), .ZN(p_wishbone_bd_ram_n25638) );
  INV_X1 U29380 ( .A(n63774), .ZN(n24910) );
  INV_X1 U29381 ( .A(n24910), .ZN(p_wishbone_bd_ram_n25637) );
  INV_X1 U29382 ( .A(n63773), .ZN(n24912) );
  INV_X1 U29383 ( .A(n24912), .ZN(p_wishbone_bd_ram_n25636) );
  INV_X1 U29384 ( .A(n63772), .ZN(n24914) );
  INV_X1 U29385 ( .A(n24914), .ZN(p_wishbone_bd_ram_n25635) );
  INV_X1 U29386 ( .A(n63771), .ZN(n24916) );
  INV_X1 U29387 ( .A(n24916), .ZN(p_wishbone_bd_ram_n25634) );
  INV_X1 U29388 ( .A(n63770), .ZN(n24918) );
  INV_X1 U29389 ( .A(n24918), .ZN(p_wishbone_bd_ram_n25633) );
  INV_X1 U29390 ( .A(n63769), .ZN(n24920) );
  INV_X1 U29391 ( .A(n24920), .ZN(p_wishbone_bd_ram_n25632) );
  INV_X1 U29392 ( .A(n63768), .ZN(n24922) );
  INV_X1 U29393 ( .A(n24922), .ZN(p_wishbone_bd_ram_n25631) );
  INV_X1 U29394 ( .A(n63767), .ZN(n24924) );
  INV_X1 U29395 ( .A(n24924), .ZN(p_wishbone_bd_ram_n25630) );
  INV_X1 U29396 ( .A(n63766), .ZN(n24926) );
  INV_X1 U29397 ( .A(n24926), .ZN(p_wishbone_bd_ram_n25629) );
  INV_X1 U29398 ( .A(n63765), .ZN(n24928) );
  INV_X1 U29399 ( .A(n24928), .ZN(p_wishbone_bd_ram_n25628) );
  INV_X1 U29400 ( .A(n63764), .ZN(n24930) );
  INV_X1 U29401 ( .A(n24930), .ZN(p_wishbone_bd_ram_n25627) );
  INV_X1 U29402 ( .A(n63763), .ZN(n24932) );
  INV_X1 U29403 ( .A(n24932), .ZN(p_wishbone_bd_ram_n25626) );
  INV_X1 U29404 ( .A(n63762), .ZN(n24934) );
  INV_X1 U29405 ( .A(n24934), .ZN(p_wishbone_bd_ram_n25625) );
  INV_X1 U29406 ( .A(n63761), .ZN(n24936) );
  INV_X1 U29407 ( .A(n24936), .ZN(p_wishbone_bd_ram_n25624) );
  INV_X1 U29408 ( .A(n63760), .ZN(n24938) );
  INV_X1 U29409 ( .A(n24938), .ZN(p_wishbone_bd_ram_n25623) );
  INV_X1 U29410 ( .A(n63759), .ZN(n24940) );
  INV_X1 U29411 ( .A(n24940), .ZN(p_wishbone_bd_ram_n25622) );
  INV_X1 U29412 ( .A(n63758), .ZN(n24942) );
  INV_X1 U29413 ( .A(n24942), .ZN(p_wishbone_bd_ram_n25621) );
  INV_X1 U29414 ( .A(n63757), .ZN(n24944) );
  INV_X1 U29415 ( .A(n24944), .ZN(p_wishbone_bd_ram_n25620) );
  INV_X1 U29416 ( .A(n63756), .ZN(n24946) );
  INV_X1 U29417 ( .A(n24946), .ZN(p_wishbone_bd_ram_n25619) );
  INV_X1 U29418 ( .A(n63755), .ZN(n24948) );
  INV_X1 U29419 ( .A(n24948), .ZN(p_wishbone_bd_ram_n25618) );
  INV_X1 U29420 ( .A(n63754), .ZN(n24950) );
  INV_X1 U29421 ( .A(n24950), .ZN(p_wishbone_bd_ram_n25617) );
  INV_X1 U29422 ( .A(n63753), .ZN(n24952) );
  INV_X1 U29423 ( .A(n24952), .ZN(p_wishbone_bd_ram_n25616) );
  INV_X1 U29424 ( .A(n63752), .ZN(n24954) );
  INV_X1 U29425 ( .A(n24954), .ZN(p_wishbone_bd_ram_n25615) );
  INV_X1 U29426 ( .A(n63751), .ZN(n24956) );
  INV_X1 U29427 ( .A(n24956), .ZN(p_wishbone_bd_ram_n25614) );
  INV_X1 U29428 ( .A(n63750), .ZN(n24958) );
  INV_X1 U29429 ( .A(n24958), .ZN(p_wishbone_bd_ram_n25613) );
  INV_X1 U29430 ( .A(n63749), .ZN(n24960) );
  INV_X1 U29431 ( .A(n24960), .ZN(p_wishbone_bd_ram_n25612) );
  INV_X1 U29432 ( .A(n63748), .ZN(n24962) );
  INV_X1 U29433 ( .A(n24962), .ZN(p_wishbone_bd_ram_n25611) );
  INV_X1 U29434 ( .A(n63747), .ZN(n24964) );
  INV_X1 U29435 ( .A(n24964), .ZN(p_wishbone_bd_ram_n25610) );
  INV_X1 U29436 ( .A(n63746), .ZN(n24966) );
  INV_X1 U29437 ( .A(n24966), .ZN(p_wishbone_bd_ram_n25609) );
  INV_X1 U29438 ( .A(n63745), .ZN(n24968) );
  INV_X1 U29439 ( .A(n24968), .ZN(p_wishbone_bd_ram_n25608) );
  INV_X1 U29440 ( .A(n63744), .ZN(n24970) );
  INV_X1 U29441 ( .A(n24970), .ZN(p_wishbone_bd_ram_n25607) );
  INV_X1 U29442 ( .A(n63743), .ZN(n24972) );
  INV_X1 U29443 ( .A(n24972), .ZN(p_wishbone_bd_ram_n25606) );
  INV_X1 U29444 ( .A(n63742), .ZN(n24974) );
  INV_X1 U29445 ( .A(n24974), .ZN(p_wishbone_bd_ram_n25605) );
  INV_X1 U29446 ( .A(n63741), .ZN(n24976) );
  INV_X1 U29447 ( .A(n24976), .ZN(p_wishbone_bd_ram_n25604) );
  INV_X1 U29448 ( .A(n63740), .ZN(n24978) );
  INV_X1 U29449 ( .A(n24978), .ZN(p_wishbone_bd_ram_n25603) );
  INV_X1 U29450 ( .A(n63739), .ZN(n24980) );
  INV_X1 U29451 ( .A(n24980), .ZN(p_wishbone_bd_ram_n25602) );
  INV_X1 U29452 ( .A(n63738), .ZN(n24982) );
  INV_X1 U29453 ( .A(n24982), .ZN(p_wishbone_bd_ram_n25601) );
  INV_X1 U29454 ( .A(n63737), .ZN(n24984) );
  INV_X1 U29455 ( .A(n24984), .ZN(p_wishbone_bd_ram_n25600) );
  INV_X1 U29456 ( .A(n63736), .ZN(n24986) );
  INV_X1 U29457 ( .A(n24986), .ZN(p_wishbone_bd_ram_n25599) );
  INV_X1 U29458 ( .A(n63735), .ZN(n24988) );
  INV_X1 U29459 ( .A(n24988), .ZN(p_wishbone_bd_ram_n25598) );
  INV_X1 U29460 ( .A(n63734), .ZN(n24990) );
  INV_X1 U29461 ( .A(n24990), .ZN(p_wishbone_bd_ram_n25597) );
  INV_X1 U29462 ( .A(n63733), .ZN(n24992) );
  INV_X1 U29463 ( .A(n24992), .ZN(p_wishbone_bd_ram_n25596) );
  INV_X1 U29464 ( .A(n63732), .ZN(n24994) );
  INV_X1 U29465 ( .A(n24994), .ZN(p_wishbone_bd_ram_n25595) );
  INV_X1 U29466 ( .A(n63731), .ZN(n24996) );
  INV_X1 U29467 ( .A(n24996), .ZN(p_wishbone_bd_ram_n25594) );
  INV_X1 U29468 ( .A(n63730), .ZN(n24998) );
  INV_X1 U29469 ( .A(n24998), .ZN(p_wishbone_bd_ram_n25593) );
  INV_X1 U29470 ( .A(n63729), .ZN(n25000) );
  INV_X1 U29471 ( .A(n25000), .ZN(p_wishbone_bd_ram_n25592) );
  INV_X1 U29472 ( .A(n63728), .ZN(n25002) );
  INV_X1 U29473 ( .A(n25002), .ZN(p_wishbone_bd_ram_n25591) );
  INV_X1 U29474 ( .A(n63727), .ZN(n25004) );
  INV_X1 U29475 ( .A(n25004), .ZN(p_wishbone_bd_ram_n25590) );
  INV_X1 U29476 ( .A(n63726), .ZN(n25006) );
  INV_X1 U29477 ( .A(n25006), .ZN(p_wishbone_bd_ram_n25589) );
  INV_X1 U29478 ( .A(n63725), .ZN(n25008) );
  INV_X1 U29479 ( .A(n25008), .ZN(p_wishbone_bd_ram_n25588) );
  INV_X1 U29480 ( .A(n63724), .ZN(n25010) );
  INV_X1 U29481 ( .A(n25010), .ZN(p_wishbone_bd_ram_n25587) );
  INV_X1 U29482 ( .A(n63723), .ZN(n25012) );
  INV_X1 U29483 ( .A(n25012), .ZN(p_wishbone_bd_ram_n25586) );
  INV_X1 U29484 ( .A(n63722), .ZN(n25014) );
  INV_X1 U29485 ( .A(n25014), .ZN(p_wishbone_bd_ram_n25585) );
  INV_X1 U29486 ( .A(n63721), .ZN(n25016) );
  INV_X1 U29487 ( .A(n25016), .ZN(p_wishbone_bd_ram_n25584) );
  INV_X1 U29488 ( .A(n63720), .ZN(n25018) );
  INV_X1 U29489 ( .A(n25018), .ZN(p_wishbone_bd_ram_n25583) );
  INV_X1 U29490 ( .A(n63719), .ZN(n25020) );
  INV_X1 U29491 ( .A(n25020), .ZN(p_wishbone_bd_ram_n25582) );
  INV_X1 U29492 ( .A(n63718), .ZN(n25022) );
  INV_X1 U29493 ( .A(n25022), .ZN(p_wishbone_bd_ram_n25581) );
  INV_X1 U29494 ( .A(n63717), .ZN(n25024) );
  INV_X1 U29495 ( .A(n25024), .ZN(p_wishbone_bd_ram_n25580) );
  INV_X1 U29496 ( .A(n63716), .ZN(n25026) );
  INV_X1 U29497 ( .A(n25026), .ZN(p_wishbone_bd_ram_n25579) );
  INV_X1 U29498 ( .A(n63715), .ZN(n25028) );
  INV_X1 U29499 ( .A(n25028), .ZN(p_wishbone_bd_ram_n25578) );
  INV_X1 U29500 ( .A(n63714), .ZN(n25030) );
  INV_X1 U29501 ( .A(n25030), .ZN(p_wishbone_bd_ram_n25577) );
  INV_X1 U29502 ( .A(n63713), .ZN(n25032) );
  INV_X1 U29503 ( .A(n25032), .ZN(p_wishbone_bd_ram_n25576) );
  INV_X1 U29504 ( .A(n63712), .ZN(n25034) );
  INV_X1 U29505 ( .A(n25034), .ZN(p_wishbone_bd_ram_n25575) );
  INV_X1 U29506 ( .A(n63711), .ZN(n25036) );
  INV_X1 U29507 ( .A(n25036), .ZN(p_wishbone_bd_ram_n25574) );
  INV_X1 U29508 ( .A(n63710), .ZN(n25038) );
  INV_X1 U29509 ( .A(n25038), .ZN(p_wishbone_bd_ram_n25573) );
  INV_X1 U29510 ( .A(n63709), .ZN(n25040) );
  INV_X1 U29511 ( .A(n25040), .ZN(p_wishbone_bd_ram_n25572) );
  INV_X1 U29512 ( .A(n63708), .ZN(n25042) );
  INV_X1 U29513 ( .A(n25042), .ZN(p_wishbone_bd_ram_n25571) );
  INV_X1 U29514 ( .A(n63707), .ZN(n25044) );
  INV_X1 U29515 ( .A(n25044), .ZN(p_wishbone_bd_ram_n25570) );
  INV_X1 U29516 ( .A(n63706), .ZN(n25046) );
  INV_X1 U29517 ( .A(n25046), .ZN(p_wishbone_bd_ram_n25569) );
  INV_X1 U29518 ( .A(n63705), .ZN(n25048) );
  INV_X1 U29519 ( .A(n25048), .ZN(p_wishbone_bd_ram_n25568) );
  INV_X1 U29520 ( .A(n63704), .ZN(n25050) );
  INV_X1 U29521 ( .A(n25050), .ZN(p_wishbone_bd_ram_n25567) );
  INV_X1 U29522 ( .A(n63703), .ZN(n25052) );
  INV_X1 U29523 ( .A(n25052), .ZN(p_wishbone_bd_ram_n25566) );
  INV_X1 U29524 ( .A(n63702), .ZN(n25054) );
  INV_X1 U29525 ( .A(n25054), .ZN(p_wishbone_bd_ram_n25565) );
  INV_X1 U29526 ( .A(n63701), .ZN(n25056) );
  INV_X1 U29527 ( .A(n25056), .ZN(p_wishbone_bd_ram_n25564) );
  INV_X1 U29528 ( .A(n63700), .ZN(n25058) );
  INV_X1 U29529 ( .A(n25058), .ZN(p_wishbone_bd_ram_n25563) );
  INV_X1 U29530 ( .A(n63699), .ZN(n25060) );
  INV_X1 U29531 ( .A(n25060), .ZN(p_wishbone_bd_ram_n25562) );
  INV_X1 U29532 ( .A(n63698), .ZN(n25062) );
  INV_X1 U29533 ( .A(n25062), .ZN(p_wishbone_bd_ram_n25561) );
  INV_X1 U29534 ( .A(n63697), .ZN(n25064) );
  INV_X1 U29535 ( .A(n25064), .ZN(p_wishbone_bd_ram_n25560) );
  INV_X1 U29536 ( .A(n63696), .ZN(n25066) );
  INV_X1 U29537 ( .A(n25066), .ZN(p_wishbone_bd_ram_n25559) );
  INV_X1 U29538 ( .A(n63695), .ZN(n25068) );
  INV_X1 U29539 ( .A(n25068), .ZN(p_wishbone_bd_ram_n25558) );
  INV_X1 U29540 ( .A(n63694), .ZN(n25070) );
  INV_X1 U29541 ( .A(n25070), .ZN(p_wishbone_bd_ram_n25557) );
  INV_X1 U29542 ( .A(n63693), .ZN(n25072) );
  INV_X1 U29543 ( .A(n25072), .ZN(p_wishbone_bd_ram_n25556) );
  INV_X1 U29544 ( .A(n63692), .ZN(n25074) );
  INV_X1 U29545 ( .A(n25074), .ZN(p_wishbone_bd_ram_n25555) );
  INV_X1 U29546 ( .A(n63691), .ZN(n25076) );
  INV_X1 U29547 ( .A(n25076), .ZN(p_wishbone_bd_ram_n25554) );
  INV_X1 U29548 ( .A(n63690), .ZN(n25078) );
  INV_X1 U29549 ( .A(n25078), .ZN(p_wishbone_bd_ram_n25553) );
  INV_X1 U29550 ( .A(n63689), .ZN(n25080) );
  INV_X1 U29551 ( .A(n25080), .ZN(p_wishbone_bd_ram_n25552) );
  INV_X1 U29552 ( .A(n63688), .ZN(n25082) );
  INV_X1 U29553 ( .A(n25082), .ZN(p_wishbone_bd_ram_n25551) );
  INV_X1 U29554 ( .A(n63687), .ZN(n25084) );
  INV_X1 U29555 ( .A(n25084), .ZN(p_wishbone_bd_ram_n25550) );
  INV_X1 U29556 ( .A(n63686), .ZN(n25086) );
  INV_X1 U29557 ( .A(n25086), .ZN(p_wishbone_bd_ram_n25549) );
  INV_X1 U29558 ( .A(n63685), .ZN(n25088) );
  INV_X1 U29559 ( .A(n25088), .ZN(p_wishbone_bd_ram_n25548) );
  INV_X1 U29560 ( .A(n63684), .ZN(n25090) );
  INV_X1 U29561 ( .A(n25090), .ZN(p_wishbone_bd_ram_n25547) );
  INV_X1 U29562 ( .A(n63683), .ZN(n25092) );
  INV_X1 U29563 ( .A(n25092), .ZN(p_wishbone_bd_ram_n25546) );
  INV_X1 U29564 ( .A(n63682), .ZN(n25094) );
  INV_X1 U29565 ( .A(n25094), .ZN(p_wishbone_bd_ram_n25545) );
  INV_X1 U29566 ( .A(n63681), .ZN(n25096) );
  INV_X1 U29567 ( .A(n25096), .ZN(p_wishbone_bd_ram_n25544) );
  INV_X1 U29568 ( .A(n63680), .ZN(n25098) );
  INV_X1 U29569 ( .A(n25098), .ZN(p_wishbone_bd_ram_n25543) );
  INV_X1 U29570 ( .A(n63679), .ZN(n25100) );
  INV_X1 U29571 ( .A(n25100), .ZN(p_wishbone_bd_ram_n25542) );
  INV_X1 U29572 ( .A(n63678), .ZN(n25102) );
  INV_X1 U29573 ( .A(n25102), .ZN(p_wishbone_bd_ram_n25541) );
  INV_X1 U29574 ( .A(n63677), .ZN(n25104) );
  INV_X1 U29575 ( .A(n25104), .ZN(p_wishbone_bd_ram_n25540) );
  INV_X1 U29576 ( .A(n63676), .ZN(n25106) );
  INV_X1 U29577 ( .A(n25106), .ZN(p_wishbone_bd_ram_n25539) );
  INV_X1 U29578 ( .A(n63675), .ZN(n25108) );
  INV_X1 U29579 ( .A(n25108), .ZN(p_wishbone_bd_ram_n25538) );
  INV_X1 U29580 ( .A(n63674), .ZN(n25110) );
  INV_X1 U29581 ( .A(n25110), .ZN(p_wishbone_bd_ram_n25537) );
  INV_X1 U29582 ( .A(n63673), .ZN(n25112) );
  INV_X1 U29583 ( .A(n25112), .ZN(p_wishbone_bd_ram_n25536) );
  INV_X1 U29584 ( .A(n63672), .ZN(n25114) );
  INV_X1 U29585 ( .A(n25114), .ZN(p_wishbone_bd_ram_n25535) );
  INV_X1 U29586 ( .A(n63671), .ZN(n25116) );
  INV_X1 U29587 ( .A(n25116), .ZN(p_wishbone_bd_ram_n25534) );
  INV_X1 U29588 ( .A(n63670), .ZN(n25118) );
  INV_X1 U29589 ( .A(n25118), .ZN(p_wishbone_bd_ram_n25533) );
  INV_X1 U29590 ( .A(n63669), .ZN(n25120) );
  INV_X1 U29591 ( .A(n25120), .ZN(p_wishbone_bd_ram_n25532) );
  INV_X1 U29592 ( .A(n63668), .ZN(n25122) );
  INV_X1 U29593 ( .A(n25122), .ZN(p_wishbone_bd_ram_n25531) );
  INV_X1 U29594 ( .A(n63667), .ZN(n25124) );
  INV_X1 U29595 ( .A(n25124), .ZN(p_wishbone_bd_ram_n25530) );
  INV_X1 U29596 ( .A(n63666), .ZN(n25126) );
  INV_X1 U29597 ( .A(n25126), .ZN(p_wishbone_bd_ram_n25529) );
  INV_X1 U29598 ( .A(n63665), .ZN(n25128) );
  INV_X1 U29599 ( .A(n25128), .ZN(p_wishbone_bd_ram_n25528) );
  INV_X1 U29600 ( .A(n63664), .ZN(n25130) );
  INV_X1 U29601 ( .A(n25130), .ZN(p_wishbone_bd_ram_n25527) );
  INV_X1 U29602 ( .A(n63663), .ZN(n25132) );
  INV_X1 U29603 ( .A(n25132), .ZN(p_wishbone_bd_ram_n25526) );
  INV_X1 U29604 ( .A(n63662), .ZN(n25134) );
  INV_X1 U29605 ( .A(n25134), .ZN(p_wishbone_bd_ram_n25525) );
  INV_X1 U29606 ( .A(n63661), .ZN(n25136) );
  INV_X1 U29607 ( .A(n25136), .ZN(p_wishbone_bd_ram_n25524) );
  INV_X1 U29608 ( .A(n63660), .ZN(n25138) );
  INV_X1 U29609 ( .A(n25138), .ZN(p_wishbone_bd_ram_n25523) );
  INV_X1 U29610 ( .A(n63659), .ZN(n25140) );
  INV_X1 U29611 ( .A(n25140), .ZN(p_wishbone_bd_ram_n25522) );
  INV_X1 U29612 ( .A(n63658), .ZN(n25142) );
  INV_X1 U29613 ( .A(n25142), .ZN(p_wishbone_bd_ram_n25521) );
  INV_X1 U29614 ( .A(n63657), .ZN(n25144) );
  INV_X1 U29615 ( .A(n25144), .ZN(p_wishbone_bd_ram_n25520) );
  INV_X1 U29616 ( .A(n63656), .ZN(n25146) );
  INV_X1 U29617 ( .A(n25146), .ZN(p_wishbone_bd_ram_n25519) );
  INV_X1 U29618 ( .A(n63655), .ZN(n25148) );
  INV_X1 U29619 ( .A(n25148), .ZN(p_wishbone_bd_ram_n25518) );
  INV_X1 U29620 ( .A(n63654), .ZN(n25150) );
  INV_X1 U29621 ( .A(n25150), .ZN(p_wishbone_bd_ram_n25517) );
  INV_X1 U29622 ( .A(n63653), .ZN(n25152) );
  INV_X1 U29623 ( .A(n25152), .ZN(p_wishbone_bd_ram_n25516) );
  INV_X1 U29624 ( .A(n63652), .ZN(n25154) );
  INV_X1 U29625 ( .A(n25154), .ZN(p_wishbone_bd_ram_n25515) );
  INV_X1 U29626 ( .A(n63651), .ZN(n25156) );
  INV_X1 U29627 ( .A(n25156), .ZN(p_wishbone_bd_ram_n25514) );
  INV_X1 U29628 ( .A(n63650), .ZN(n25158) );
  INV_X1 U29629 ( .A(n25158), .ZN(p_wishbone_bd_ram_n25513) );
  INV_X1 U29630 ( .A(n63649), .ZN(n25160) );
  INV_X1 U29631 ( .A(n25160), .ZN(p_wishbone_bd_ram_n25512) );
  INV_X1 U29632 ( .A(n63648), .ZN(n25162) );
  INV_X1 U29633 ( .A(n25162), .ZN(p_wishbone_bd_ram_n25511) );
  INV_X1 U29634 ( .A(n63647), .ZN(n25164) );
  INV_X1 U29635 ( .A(n25164), .ZN(p_wishbone_bd_ram_n25510) );
  INV_X1 U29636 ( .A(n63646), .ZN(n25166) );
  INV_X1 U29637 ( .A(n25166), .ZN(p_wishbone_bd_ram_n25509) );
  INV_X1 U29638 ( .A(n63645), .ZN(n25168) );
  INV_X1 U29639 ( .A(n25168), .ZN(p_wishbone_bd_ram_n25508) );
  INV_X1 U29640 ( .A(n63644), .ZN(n25170) );
  INV_X1 U29641 ( .A(n25170), .ZN(p_wishbone_bd_ram_n25507) );
  INV_X1 U29642 ( .A(n63643), .ZN(n25172) );
  INV_X1 U29643 ( .A(n25172), .ZN(p_wishbone_bd_ram_n25506) );
  INV_X1 U29644 ( .A(n63642), .ZN(n25174) );
  INV_X1 U29645 ( .A(n25174), .ZN(p_wishbone_bd_ram_n25505) );
  INV_X1 U29646 ( .A(n63641), .ZN(n25176) );
  INV_X1 U29647 ( .A(n25176), .ZN(p_wishbone_bd_ram_n25504) );
  INV_X1 U29648 ( .A(n63640), .ZN(n25178) );
  INV_X1 U29649 ( .A(n25178), .ZN(p_wishbone_bd_ram_n25503) );
  INV_X1 U29650 ( .A(n63639), .ZN(n25180) );
  INV_X1 U29651 ( .A(n25180), .ZN(p_wishbone_bd_ram_n25502) );
  INV_X1 U29652 ( .A(n63638), .ZN(n25182) );
  INV_X1 U29653 ( .A(n25182), .ZN(p_wishbone_bd_ram_n25501) );
  INV_X1 U29654 ( .A(n63637), .ZN(n25184) );
  INV_X1 U29655 ( .A(n25184), .ZN(p_wishbone_bd_ram_n25500) );
  INV_X1 U29656 ( .A(n63636), .ZN(n25186) );
  INV_X1 U29657 ( .A(n25186), .ZN(p_wishbone_bd_ram_n25499) );
  INV_X1 U29658 ( .A(n63635), .ZN(n25188) );
  INV_X1 U29659 ( .A(n25188), .ZN(p_wishbone_bd_ram_n25498) );
  INV_X1 U29660 ( .A(n63634), .ZN(n25190) );
  INV_X1 U29661 ( .A(n25190), .ZN(p_wishbone_bd_ram_n25497) );
  INV_X1 U29662 ( .A(n63633), .ZN(n25192) );
  INV_X1 U29663 ( .A(n25192), .ZN(p_wishbone_bd_ram_n25496) );
  INV_X1 U29664 ( .A(n63632), .ZN(n25194) );
  INV_X1 U29665 ( .A(n25194), .ZN(p_wishbone_bd_ram_n25495) );
  INV_X1 U29666 ( .A(n63631), .ZN(n25196) );
  INV_X1 U29667 ( .A(n25196), .ZN(p_wishbone_bd_ram_n25494) );
  INV_X1 U29668 ( .A(n63630), .ZN(n25198) );
  INV_X1 U29669 ( .A(n25198), .ZN(p_wishbone_bd_ram_n25493) );
  INV_X1 U29670 ( .A(n63629), .ZN(n25200) );
  INV_X1 U29671 ( .A(n25200), .ZN(p_wishbone_bd_ram_n25492) );
  INV_X1 U29672 ( .A(n63628), .ZN(n25202) );
  INV_X1 U29673 ( .A(n25202), .ZN(p_wishbone_bd_ram_n25491) );
  INV_X1 U29674 ( .A(n63627), .ZN(n25204) );
  INV_X1 U29675 ( .A(n25204), .ZN(p_wishbone_bd_ram_n25490) );
  INV_X1 U29676 ( .A(n63626), .ZN(n25206) );
  INV_X1 U29677 ( .A(n25206), .ZN(p_wishbone_bd_ram_n25489) );
  INV_X1 U29678 ( .A(n63625), .ZN(n25208) );
  INV_X1 U29679 ( .A(n25208), .ZN(p_wishbone_bd_ram_n25488) );
  INV_X1 U29680 ( .A(n63624), .ZN(n25210) );
  INV_X1 U29681 ( .A(n25210), .ZN(p_wishbone_bd_ram_n25487) );
  INV_X1 U29682 ( .A(n63623), .ZN(n25212) );
  INV_X1 U29683 ( .A(n25212), .ZN(p_wishbone_bd_ram_n25486) );
  INV_X1 U29684 ( .A(n63622), .ZN(n25214) );
  INV_X1 U29685 ( .A(n25214), .ZN(p_wishbone_bd_ram_n25485) );
  INV_X1 U29686 ( .A(n63621), .ZN(n25216) );
  INV_X1 U29687 ( .A(n25216), .ZN(p_wishbone_bd_ram_n25484) );
  INV_X1 U29688 ( .A(n63620), .ZN(n25218) );
  INV_X1 U29689 ( .A(n25218), .ZN(p_wishbone_bd_ram_n25483) );
  INV_X1 U29690 ( .A(n63619), .ZN(n25220) );
  INV_X1 U29691 ( .A(n25220), .ZN(p_wishbone_bd_ram_n25482) );
  INV_X1 U29692 ( .A(n63618), .ZN(n25222) );
  INV_X1 U29693 ( .A(n25222), .ZN(p_wishbone_bd_ram_n25481) );
  INV_X1 U29694 ( .A(n63617), .ZN(n25224) );
  INV_X1 U29695 ( .A(n25224), .ZN(p_wishbone_bd_ram_n25480) );
  INV_X1 U29696 ( .A(n63616), .ZN(n25226) );
  INV_X1 U29697 ( .A(n25226), .ZN(p_wishbone_bd_ram_n25479) );
  INV_X1 U29698 ( .A(n63615), .ZN(n25228) );
  INV_X1 U29699 ( .A(n25228), .ZN(p_wishbone_bd_ram_n25478) );
  INV_X1 U29700 ( .A(n63614), .ZN(n25230) );
  INV_X1 U29701 ( .A(n25230), .ZN(p_wishbone_bd_ram_n25477) );
  INV_X1 U29702 ( .A(n63613), .ZN(n25232) );
  INV_X1 U29703 ( .A(n25232), .ZN(p_wishbone_bd_ram_n25476) );
  INV_X1 U29704 ( .A(n63612), .ZN(n25234) );
  INV_X1 U29705 ( .A(n25234), .ZN(p_wishbone_bd_ram_n25475) );
  INV_X1 U29706 ( .A(n63611), .ZN(n25236) );
  INV_X1 U29707 ( .A(n25236), .ZN(p_wishbone_bd_ram_n25474) );
  INV_X1 U29708 ( .A(n63610), .ZN(n25238) );
  INV_X1 U29709 ( .A(n25238), .ZN(p_wishbone_bd_ram_n25473) );
  INV_X1 U29710 ( .A(n63609), .ZN(n25240) );
  INV_X1 U29711 ( .A(n25240), .ZN(p_wishbone_bd_ram_n25472) );
  INV_X1 U29712 ( .A(n63608), .ZN(n25242) );
  INV_X1 U29713 ( .A(n25242), .ZN(p_wishbone_bd_ram_n25471) );
  INV_X1 U29714 ( .A(n63607), .ZN(n25244) );
  INV_X1 U29715 ( .A(n25244), .ZN(p_wishbone_bd_ram_n25470) );
  INV_X1 U29716 ( .A(n63606), .ZN(n25246) );
  INV_X1 U29717 ( .A(n25246), .ZN(p_wishbone_bd_ram_n25469) );
  INV_X1 U29718 ( .A(n63605), .ZN(n25248) );
  INV_X1 U29719 ( .A(n25248), .ZN(p_wishbone_bd_ram_n25468) );
  INV_X1 U29720 ( .A(n63604), .ZN(n25250) );
  INV_X1 U29721 ( .A(n25250), .ZN(p_wishbone_bd_ram_n25467) );
  INV_X1 U29722 ( .A(n63603), .ZN(n25252) );
  INV_X1 U29723 ( .A(n25252), .ZN(p_wishbone_bd_ram_n25466) );
  INV_X1 U29724 ( .A(n63602), .ZN(n25254) );
  INV_X1 U29725 ( .A(n25254), .ZN(p_wishbone_bd_ram_n25465) );
  INV_X1 U29726 ( .A(n63601), .ZN(n25256) );
  INV_X1 U29727 ( .A(n25256), .ZN(p_wishbone_bd_ram_n25464) );
  INV_X1 U29728 ( .A(n63600), .ZN(n25258) );
  INV_X1 U29729 ( .A(n25258), .ZN(p_wishbone_bd_ram_n25463) );
  INV_X1 U29730 ( .A(n63599), .ZN(n25260) );
  INV_X1 U29731 ( .A(n25260), .ZN(p_wishbone_bd_ram_n25462) );
  INV_X1 U29732 ( .A(n63598), .ZN(n25262) );
  INV_X1 U29733 ( .A(n25262), .ZN(p_wishbone_bd_ram_n25461) );
  INV_X1 U29734 ( .A(n63597), .ZN(n25264) );
  INV_X1 U29735 ( .A(n25264), .ZN(p_wishbone_bd_ram_n25460) );
  INV_X1 U29736 ( .A(n63596), .ZN(n25266) );
  INV_X1 U29737 ( .A(n25266), .ZN(p_wishbone_bd_ram_n25459) );
  INV_X1 U29738 ( .A(n63595), .ZN(n25268) );
  INV_X1 U29739 ( .A(n25268), .ZN(p_wishbone_bd_ram_n25458) );
  INV_X1 U29740 ( .A(n63594), .ZN(n25270) );
  INV_X1 U29741 ( .A(n25270), .ZN(p_wishbone_bd_ram_n25457) );
  INV_X1 U29742 ( .A(n63593), .ZN(n25272) );
  INV_X1 U29743 ( .A(n25272), .ZN(p_wishbone_bd_ram_n25456) );
  INV_X1 U29744 ( .A(n63592), .ZN(n25274) );
  INV_X1 U29745 ( .A(n25274), .ZN(p_wishbone_bd_ram_n25455) );
  INV_X1 U29746 ( .A(n63591), .ZN(n25276) );
  INV_X1 U29747 ( .A(n25276), .ZN(p_wishbone_bd_ram_n25454) );
  INV_X1 U29748 ( .A(n63590), .ZN(n25278) );
  INV_X1 U29749 ( .A(n25278), .ZN(p_wishbone_bd_ram_n25453) );
  INV_X1 U29750 ( .A(n63589), .ZN(n25280) );
  INV_X1 U29751 ( .A(n25280), .ZN(p_wishbone_bd_ram_n25452) );
  INV_X1 U29752 ( .A(n63588), .ZN(n25282) );
  INV_X1 U29753 ( .A(n25282), .ZN(p_wishbone_bd_ram_n25451) );
  INV_X1 U29754 ( .A(n63587), .ZN(n25284) );
  INV_X1 U29755 ( .A(n25284), .ZN(p_wishbone_bd_ram_n25450) );
  INV_X1 U29756 ( .A(n63586), .ZN(n25286) );
  INV_X1 U29757 ( .A(n25286), .ZN(p_wishbone_bd_ram_n25449) );
  INV_X1 U29758 ( .A(n63585), .ZN(n25288) );
  INV_X1 U29759 ( .A(n25288), .ZN(p_wishbone_bd_ram_n25448) );
  INV_X1 U29760 ( .A(n63584), .ZN(n25290) );
  INV_X1 U29761 ( .A(n25290), .ZN(p_wishbone_bd_ram_n25447) );
  INV_X1 U29762 ( .A(n63583), .ZN(n25292) );
  INV_X1 U29763 ( .A(n25292), .ZN(p_wishbone_bd_ram_n25446) );
  INV_X1 U29764 ( .A(n63582), .ZN(n25294) );
  INV_X1 U29765 ( .A(n25294), .ZN(p_wishbone_bd_ram_n25445) );
  INV_X1 U29766 ( .A(n63581), .ZN(n25296) );
  INV_X1 U29767 ( .A(n25296), .ZN(p_wishbone_bd_ram_n25444) );
  INV_X1 U29768 ( .A(n63580), .ZN(n25298) );
  INV_X1 U29769 ( .A(n25298), .ZN(p_wishbone_bd_ram_n25443) );
  INV_X1 U29770 ( .A(n63579), .ZN(n25300) );
  INV_X1 U29771 ( .A(n25300), .ZN(p_wishbone_bd_ram_n25442) );
  INV_X1 U29772 ( .A(n63578), .ZN(n25302) );
  INV_X1 U29773 ( .A(n25302), .ZN(p_wishbone_bd_ram_n25441) );
  INV_X1 U29774 ( .A(n63577), .ZN(n25304) );
  INV_X1 U29775 ( .A(n25304), .ZN(p_wishbone_bd_ram_n25440) );
  INV_X1 U29776 ( .A(n63576), .ZN(n25306) );
  INV_X1 U29777 ( .A(n25306), .ZN(p_wishbone_bd_ram_n25439) );
  INV_X1 U29778 ( .A(n63575), .ZN(n25308) );
  INV_X1 U29779 ( .A(n25308), .ZN(p_wishbone_bd_ram_n25438) );
  INV_X1 U29780 ( .A(n63574), .ZN(n25310) );
  INV_X1 U29781 ( .A(n25310), .ZN(p_wishbone_bd_ram_n25437) );
  INV_X1 U29782 ( .A(n63573), .ZN(n25312) );
  INV_X1 U29783 ( .A(n25312), .ZN(p_wishbone_bd_ram_n25436) );
  INV_X1 U29784 ( .A(n63572), .ZN(n25314) );
  INV_X1 U29785 ( .A(n25314), .ZN(p_wishbone_bd_ram_n25435) );
  INV_X1 U29786 ( .A(n63571), .ZN(n25316) );
  INV_X1 U29787 ( .A(n25316), .ZN(p_wishbone_bd_ram_n25434) );
  INV_X1 U29788 ( .A(n63570), .ZN(n25318) );
  INV_X1 U29789 ( .A(n25318), .ZN(p_wishbone_bd_ram_n25433) );
  INV_X1 U29790 ( .A(n63569), .ZN(n25320) );
  INV_X1 U29791 ( .A(n25320), .ZN(p_wishbone_bd_ram_n25432) );
  INV_X1 U29792 ( .A(n63568), .ZN(n25322) );
  INV_X1 U29793 ( .A(n25322), .ZN(p_wishbone_bd_ram_n25431) );
  INV_X1 U29794 ( .A(n63567), .ZN(n25324) );
  INV_X1 U29795 ( .A(n25324), .ZN(p_wishbone_bd_ram_n25430) );
  INV_X1 U29796 ( .A(n63566), .ZN(n25326) );
  INV_X1 U29797 ( .A(n25326), .ZN(p_wishbone_bd_ram_n25429) );
  INV_X1 U29798 ( .A(n63565), .ZN(n25328) );
  INV_X1 U29799 ( .A(n25328), .ZN(p_wishbone_bd_ram_n25428) );
  INV_X1 U29800 ( .A(n63564), .ZN(n25330) );
  INV_X1 U29801 ( .A(n25330), .ZN(p_wishbone_bd_ram_n25427) );
  INV_X1 U29802 ( .A(n63563), .ZN(n25332) );
  INV_X1 U29803 ( .A(n25332), .ZN(p_wishbone_bd_ram_n25426) );
  INV_X1 U29804 ( .A(n63562), .ZN(n25334) );
  INV_X1 U29805 ( .A(n25334), .ZN(p_wishbone_bd_ram_n25425) );
  INV_X1 U29806 ( .A(n63561), .ZN(n25336) );
  INV_X1 U29807 ( .A(n25336), .ZN(p_wishbone_bd_ram_n25424) );
  INV_X1 U29808 ( .A(n63560), .ZN(n25338) );
  INV_X1 U29809 ( .A(n25338), .ZN(p_wishbone_bd_ram_n25423) );
  INV_X1 U29810 ( .A(n63559), .ZN(n25340) );
  INV_X1 U29811 ( .A(n25340), .ZN(p_wishbone_bd_ram_n25422) );
  INV_X1 U29812 ( .A(n63558), .ZN(n25342) );
  INV_X1 U29813 ( .A(n25342), .ZN(p_wishbone_bd_ram_n25421) );
  INV_X1 U29814 ( .A(n63557), .ZN(n25344) );
  INV_X1 U29815 ( .A(n25344), .ZN(p_wishbone_bd_ram_n25420) );
  INV_X1 U29816 ( .A(n63556), .ZN(n25346) );
  INV_X1 U29817 ( .A(n25346), .ZN(p_wishbone_bd_ram_n25419) );
  INV_X1 U29818 ( .A(n63555), .ZN(n25348) );
  INV_X1 U29819 ( .A(n25348), .ZN(p_wishbone_bd_ram_n25418) );
  INV_X1 U29820 ( .A(n63554), .ZN(n25350) );
  INV_X1 U29821 ( .A(n25350), .ZN(p_wishbone_bd_ram_n25417) );
  INV_X1 U29822 ( .A(n63553), .ZN(n25352) );
  INV_X1 U29823 ( .A(n25352), .ZN(p_wishbone_bd_ram_n25416) );
  INV_X1 U29824 ( .A(n63552), .ZN(n25354) );
  INV_X1 U29825 ( .A(n25354), .ZN(p_wishbone_bd_ram_n25415) );
  INV_X1 U29826 ( .A(n63551), .ZN(n25356) );
  INV_X1 U29827 ( .A(n25356), .ZN(p_wishbone_bd_ram_n25414) );
  INV_X1 U29828 ( .A(n63550), .ZN(n25358) );
  INV_X1 U29829 ( .A(n25358), .ZN(p_wishbone_bd_ram_n25413) );
  INV_X1 U29830 ( .A(n63549), .ZN(n25360) );
  INV_X1 U29831 ( .A(n25360), .ZN(p_wishbone_bd_ram_n25412) );
  INV_X1 U29832 ( .A(n63548), .ZN(n25362) );
  INV_X1 U29833 ( .A(n25362), .ZN(p_wishbone_bd_ram_n25411) );
  INV_X1 U29834 ( .A(n63547), .ZN(n25364) );
  INV_X1 U29835 ( .A(n25364), .ZN(p_wishbone_bd_ram_n25410) );
  INV_X1 U29836 ( .A(n63546), .ZN(n25366) );
  INV_X1 U29837 ( .A(n25366), .ZN(p_wishbone_bd_ram_n25409) );
  INV_X1 U29838 ( .A(n63545), .ZN(n25368) );
  INV_X1 U29839 ( .A(n25368), .ZN(p_wishbone_bd_ram_n25408) );
  INV_X1 U29840 ( .A(n63544), .ZN(n25370) );
  INV_X1 U29841 ( .A(n25370), .ZN(p_wishbone_bd_ram_n25407) );
  INV_X1 U29842 ( .A(n63543), .ZN(n25372) );
  INV_X1 U29843 ( .A(n25372), .ZN(p_wishbone_bd_ram_n25406) );
  INV_X1 U29844 ( .A(n63542), .ZN(n25374) );
  INV_X1 U29845 ( .A(n25374), .ZN(p_wishbone_bd_ram_n25405) );
  INV_X1 U29846 ( .A(n63541), .ZN(n25376) );
  INV_X1 U29847 ( .A(n25376), .ZN(p_wishbone_bd_ram_n25404) );
  INV_X1 U29848 ( .A(n63540), .ZN(n25378) );
  INV_X1 U29849 ( .A(n25378), .ZN(p_wishbone_bd_ram_n25403) );
  INV_X1 U29850 ( .A(n63539), .ZN(n25380) );
  INV_X1 U29851 ( .A(n25380), .ZN(p_wishbone_bd_ram_n25402) );
  INV_X1 U29852 ( .A(n63538), .ZN(n25382) );
  INV_X1 U29853 ( .A(n25382), .ZN(p_wishbone_bd_ram_n25401) );
  INV_X1 U29854 ( .A(n63537), .ZN(n25384) );
  INV_X1 U29855 ( .A(n25384), .ZN(p_wishbone_bd_ram_n25400) );
  INV_X1 U29856 ( .A(n63536), .ZN(n25386) );
  INV_X1 U29857 ( .A(n25386), .ZN(p_wishbone_bd_ram_n25399) );
  INV_X1 U29858 ( .A(n63535), .ZN(n25388) );
  INV_X1 U29859 ( .A(n25388), .ZN(p_wishbone_bd_ram_n25398) );
  INV_X1 U29860 ( .A(n63534), .ZN(n25390) );
  INV_X1 U29861 ( .A(n25390), .ZN(p_wishbone_bd_ram_n25397) );
  INV_X1 U29862 ( .A(n63533), .ZN(n25392) );
  INV_X1 U29863 ( .A(n25392), .ZN(p_wishbone_bd_ram_n25396) );
  INV_X1 U29864 ( .A(n63532), .ZN(n25394) );
  INV_X1 U29865 ( .A(n25394), .ZN(p_wishbone_bd_ram_n25395) );
  INV_X1 U29866 ( .A(n63531), .ZN(n25396) );
  INV_X1 U29867 ( .A(n25396), .ZN(p_wishbone_bd_ram_n25394) );
  INV_X1 U29868 ( .A(n63530), .ZN(n25398) );
  INV_X1 U29869 ( .A(n25398), .ZN(p_wishbone_bd_ram_n25393) );
  INV_X1 U29870 ( .A(n63529), .ZN(n25400) );
  INV_X1 U29871 ( .A(n25400), .ZN(p_wishbone_bd_ram_n25392) );
  INV_X1 U29872 ( .A(n63528), .ZN(n25402) );
  INV_X1 U29873 ( .A(n25402), .ZN(p_wishbone_bd_ram_n25391) );
  INV_X1 U29874 ( .A(n63527), .ZN(n25404) );
  INV_X1 U29875 ( .A(n25404), .ZN(p_wishbone_bd_ram_n25390) );
  INV_X1 U29876 ( .A(n63526), .ZN(n25406) );
  INV_X1 U29877 ( .A(n25406), .ZN(p_wishbone_bd_ram_n25389) );
  INV_X1 U29878 ( .A(n63525), .ZN(n25408) );
  INV_X1 U29879 ( .A(n25408), .ZN(p_wishbone_bd_ram_n25388) );
  INV_X1 U29880 ( .A(n63524), .ZN(n25410) );
  INV_X1 U29881 ( .A(n25410), .ZN(p_wishbone_bd_ram_n25387) );
  INV_X1 U29882 ( .A(n63523), .ZN(n25412) );
  INV_X1 U29883 ( .A(n25412), .ZN(p_wishbone_bd_ram_n25386) );
  INV_X1 U29884 ( .A(n63522), .ZN(n25414) );
  INV_X1 U29885 ( .A(n25414), .ZN(p_wishbone_bd_ram_n25385) );
  INV_X1 U29886 ( .A(n63521), .ZN(n25416) );
  INV_X1 U29887 ( .A(n25416), .ZN(p_wishbone_bd_ram_n25384) );
  INV_X1 U29888 ( .A(n63520), .ZN(n25418) );
  INV_X1 U29889 ( .A(n25418), .ZN(p_wishbone_bd_ram_n25383) );
  INV_X1 U29890 ( .A(n63519), .ZN(n25420) );
  INV_X1 U29891 ( .A(n25420), .ZN(p_wishbone_bd_ram_n25382) );
  INV_X1 U29892 ( .A(n63518), .ZN(n25422) );
  INV_X1 U29893 ( .A(n25422), .ZN(p_wishbone_bd_ram_n25381) );
  INV_X1 U29894 ( .A(n63517), .ZN(n25424) );
  INV_X1 U29895 ( .A(n25424), .ZN(p_wishbone_bd_ram_n25380) );
  INV_X1 U29896 ( .A(n63516), .ZN(n25426) );
  INV_X1 U29897 ( .A(n25426), .ZN(p_wishbone_bd_ram_n25379) );
  INV_X1 U29898 ( .A(n63515), .ZN(n25428) );
  INV_X1 U29899 ( .A(n25428), .ZN(p_wishbone_bd_ram_n25378) );
  INV_X1 U29900 ( .A(n63514), .ZN(n25430) );
  INV_X1 U29901 ( .A(n25430), .ZN(p_wishbone_bd_ram_n25377) );
  INV_X1 U29902 ( .A(n63513), .ZN(n25432) );
  INV_X1 U29903 ( .A(n25432), .ZN(p_wishbone_bd_ram_n25376) );
  INV_X1 U29904 ( .A(n63512), .ZN(n25434) );
  INV_X1 U29905 ( .A(n25434), .ZN(p_wishbone_bd_ram_n25375) );
  INV_X1 U29906 ( .A(n63511), .ZN(n25436) );
  INV_X1 U29907 ( .A(n25436), .ZN(p_wishbone_bd_ram_n25374) );
  INV_X1 U29908 ( .A(n63510), .ZN(n25438) );
  INV_X1 U29909 ( .A(n25438), .ZN(p_wishbone_bd_ram_n25373) );
  INV_X1 U29910 ( .A(n63509), .ZN(n25440) );
  INV_X1 U29911 ( .A(n25440), .ZN(p_wishbone_bd_ram_n25372) );
  INV_X1 U29912 ( .A(n63508), .ZN(n25442) );
  INV_X1 U29913 ( .A(n25442), .ZN(p_wishbone_bd_ram_n25371) );
  INV_X1 U29914 ( .A(n63507), .ZN(n25444) );
  INV_X1 U29915 ( .A(n25444), .ZN(p_wishbone_bd_ram_n25370) );
  INV_X1 U29916 ( .A(n63506), .ZN(n25446) );
  INV_X1 U29917 ( .A(n25446), .ZN(p_wishbone_bd_ram_n25369) );
  INV_X1 U29918 ( .A(n63505), .ZN(n25448) );
  INV_X1 U29919 ( .A(n25448), .ZN(p_wishbone_bd_ram_n25368) );
  INV_X1 U29920 ( .A(n63504), .ZN(n25450) );
  INV_X1 U29921 ( .A(n25450), .ZN(p_wishbone_bd_ram_n25367) );
  INV_X1 U29922 ( .A(n63503), .ZN(n25452) );
  INV_X1 U29923 ( .A(n25452), .ZN(p_wishbone_bd_ram_n25366) );
  INV_X1 U29924 ( .A(n63502), .ZN(n25454) );
  INV_X1 U29925 ( .A(n25454), .ZN(p_wishbone_bd_ram_n25365) );
  INV_X1 U29926 ( .A(n63501), .ZN(n25456) );
  INV_X1 U29927 ( .A(n25456), .ZN(p_wishbone_bd_ram_n25364) );
  INV_X1 U29928 ( .A(n63500), .ZN(n25458) );
  INV_X1 U29929 ( .A(n25458), .ZN(p_wishbone_bd_ram_n25363) );
  INV_X1 U29930 ( .A(n63499), .ZN(n25460) );
  INV_X1 U29931 ( .A(n25460), .ZN(p_wishbone_bd_ram_n25362) );
  INV_X1 U29932 ( .A(n63498), .ZN(n25462) );
  INV_X1 U29933 ( .A(n25462), .ZN(p_wishbone_bd_ram_n25361) );
  INV_X1 U29934 ( .A(n63497), .ZN(n25464) );
  INV_X1 U29935 ( .A(n25464), .ZN(p_wishbone_bd_ram_n25359) );
  INV_X1 U29936 ( .A(n63496), .ZN(n25466) );
  INV_X1 U29937 ( .A(n25466), .ZN(p_wishbone_bd_ram_n25357) );
  INV_X1 U29938 ( .A(n63495), .ZN(n25468) );
  INV_X1 U29939 ( .A(n25468), .ZN(p_wishbone_bd_ram_n25356) );
  INV_X1 U29940 ( .A(n63494), .ZN(n25470) );
  INV_X1 U29941 ( .A(n25470), .ZN(p_wishbone_bd_ram_n25354) );
  INV_X1 U29942 ( .A(n63493), .ZN(n25472) );
  INV_X1 U29943 ( .A(n25472), .ZN(p_wishbone_bd_ram_n25352) );
  INV_X1 U29944 ( .A(n63492), .ZN(n25474) );
  INV_X1 U29945 ( .A(n25474), .ZN(p_wishbone_bd_ram_n25351) );
  INV_X1 U29946 ( .A(n63491), .ZN(n25476) );
  INV_X1 U29947 ( .A(n25476), .ZN(p_wishbone_bd_ram_n25350) );
  INV_X1 U29948 ( .A(n63490), .ZN(n25478) );
  INV_X1 U29949 ( .A(n25478), .ZN(p_wishbone_bd_ram_n25349) );
  INV_X1 U29950 ( .A(n63489), .ZN(n25480) );
  INV_X1 U29951 ( .A(n25480), .ZN(p_wishbone_bd_ram_n25348) );
  INV_X1 U29952 ( .A(n63488), .ZN(n25482) );
  INV_X1 U29953 ( .A(n25482), .ZN(p_wishbone_bd_ram_n25347) );
  INV_X1 U29954 ( .A(n63487), .ZN(n25484) );
  INV_X1 U29955 ( .A(n25484), .ZN(p_wishbone_bd_ram_n25346) );
  INV_X1 U29956 ( .A(n63486), .ZN(n25486) );
  INV_X1 U29957 ( .A(n25486), .ZN(p_wishbone_bd_ram_n25345) );
  INV_X1 U29958 ( .A(n63485), .ZN(n25488) );
  INV_X1 U29959 ( .A(n25488), .ZN(p_wishbone_bd_ram_n25344) );
  INV_X1 U29960 ( .A(n63484), .ZN(n25490) );
  INV_X1 U29961 ( .A(n25490), .ZN(p_wishbone_bd_ram_n25343) );
  INV_X1 U29962 ( .A(n63483), .ZN(n25492) );
  INV_X1 U29963 ( .A(n25492), .ZN(p_wishbone_bd_ram_n25342) );
  INV_X1 U29964 ( .A(n63482), .ZN(n25494) );
  INV_X1 U29965 ( .A(n25494), .ZN(p_wishbone_bd_ram_n25341) );
  INV_X1 U29966 ( .A(n63481), .ZN(n25496) );
  INV_X1 U29967 ( .A(n25496), .ZN(p_wishbone_bd_ram_n25340) );
  INV_X1 U29968 ( .A(n63480), .ZN(n25498) );
  INV_X1 U29969 ( .A(n25498), .ZN(p_wishbone_bd_ram_n25339) );
  INV_X1 U29970 ( .A(n63479), .ZN(n25500) );
  INV_X1 U29971 ( .A(n25500), .ZN(p_wishbone_bd_ram_n25338) );
  INV_X1 U29972 ( .A(n63478), .ZN(n25502) );
  INV_X1 U29973 ( .A(n25502), .ZN(p_wishbone_bd_ram_n25337) );
  INV_X1 U29974 ( .A(n63477), .ZN(n25504) );
  INV_X1 U29975 ( .A(n25504), .ZN(p_wishbone_bd_ram_n25336) );
  INV_X1 U29976 ( .A(n63476), .ZN(n25506) );
  INV_X1 U29977 ( .A(n25506), .ZN(p_wishbone_bd_ram_n25335) );
  INV_X1 U29978 ( .A(n63475), .ZN(n25508) );
  INV_X1 U29979 ( .A(n25508), .ZN(p_wishbone_bd_ram_n25334) );
  INV_X1 U29980 ( .A(n63474), .ZN(n25510) );
  INV_X1 U29981 ( .A(n25510), .ZN(p_wishbone_bd_ram_n25333) );
  INV_X1 U29982 ( .A(n63473), .ZN(n25512) );
  INV_X1 U29983 ( .A(n25512), .ZN(p_wishbone_bd_ram_n25332) );
  INV_X1 U29984 ( .A(n63472), .ZN(n25514) );
  INV_X1 U29985 ( .A(n25514), .ZN(p_wishbone_bd_ram_n25331) );
  INV_X1 U29986 ( .A(n63471), .ZN(n25516) );
  INV_X1 U29987 ( .A(n25516), .ZN(p_wishbone_bd_ram_n25330) );
  INV_X1 U29988 ( .A(n63470), .ZN(n25518) );
  INV_X1 U29989 ( .A(n25518), .ZN(p_wishbone_bd_ram_n25329) );
  INV_X1 U29990 ( .A(n63469), .ZN(n25520) );
  INV_X1 U29991 ( .A(n25520), .ZN(p_wishbone_bd_ram_n25328) );
  INV_X1 U29992 ( .A(n63468), .ZN(n25522) );
  INV_X1 U29993 ( .A(n25522), .ZN(p_wishbone_bd_ram_n25327) );
  INV_X1 U29994 ( .A(n63467), .ZN(n25524) );
  INV_X1 U29995 ( .A(n25524), .ZN(p_wishbone_bd_ram_n25326) );
  INV_X1 U29996 ( .A(n63466), .ZN(n25526) );
  INV_X1 U29997 ( .A(n25526), .ZN(p_wishbone_bd_ram_n25325) );
  INV_X1 U29998 ( .A(n63465), .ZN(n25528) );
  INV_X1 U29999 ( .A(n25528), .ZN(p_wishbone_bd_ram_n25324) );
  INV_X1 U30000 ( .A(n63464), .ZN(n25530) );
  INV_X1 U30001 ( .A(n25530), .ZN(p_wishbone_bd_ram_n25323) );
  INV_X1 U30002 ( .A(n63463), .ZN(n25532) );
  INV_X1 U30003 ( .A(n25532), .ZN(p_wishbone_bd_ram_n25322) );
  INV_X1 U30004 ( .A(n63462), .ZN(n25534) );
  INV_X1 U30005 ( .A(n25534), .ZN(p_wishbone_bd_ram_n25321) );
  INV_X1 U30006 ( .A(n63461), .ZN(n25536) );
  INV_X1 U30007 ( .A(n25536), .ZN(p_wishbone_bd_ram_n25320) );
  INV_X1 U30008 ( .A(n63460), .ZN(n25538) );
  INV_X1 U30009 ( .A(n25538), .ZN(p_wishbone_bd_ram_n25319) );
  INV_X1 U30010 ( .A(n63459), .ZN(n25540) );
  INV_X1 U30011 ( .A(n25540), .ZN(p_wishbone_bd_ram_n25318) );
  INV_X1 U30012 ( .A(n63458), .ZN(n25542) );
  INV_X1 U30013 ( .A(n25542), .ZN(p_wishbone_bd_ram_n25317) );
  INV_X1 U30014 ( .A(n63457), .ZN(n25544) );
  INV_X1 U30015 ( .A(n25544), .ZN(p_wishbone_bd_ram_n25316) );
  INV_X1 U30016 ( .A(n63456), .ZN(n25546) );
  INV_X1 U30017 ( .A(n25546), .ZN(p_wishbone_bd_ram_n25315) );
  INV_X1 U30018 ( .A(n63455), .ZN(n25548) );
  INV_X1 U30019 ( .A(n25548), .ZN(p_wishbone_bd_ram_n25314) );
  INV_X1 U30020 ( .A(n63454), .ZN(n25550) );
  INV_X1 U30021 ( .A(n25550), .ZN(p_wishbone_bd_ram_n25313) );
  INV_X1 U30022 ( .A(n63453), .ZN(n25552) );
  INV_X1 U30023 ( .A(n25552), .ZN(p_wishbone_bd_ram_n25312) );
  INV_X1 U30024 ( .A(n63452), .ZN(n25554) );
  INV_X1 U30025 ( .A(n25554), .ZN(p_wishbone_bd_ram_n25310) );
  INV_X1 U30026 ( .A(n63451), .ZN(n25556) );
  INV_X1 U30027 ( .A(n25556), .ZN(p_wishbone_bd_ram_n25307) );
  INV_X1 U30028 ( .A(n63450), .ZN(n25558) );
  INV_X1 U30029 ( .A(n25558), .ZN(p_wishbone_bd_ram_n25305) );
  INV_X1 U30030 ( .A(n63449), .ZN(n25560) );
  INV_X1 U30031 ( .A(n25560), .ZN(p_wishbone_bd_ram_n25304) );
  INV_X1 U30032 ( .A(n63448), .ZN(n25562) );
  INV_X1 U30033 ( .A(n25562), .ZN(p_wishbone_bd_ram_n25303) );
  INV_X1 U30034 ( .A(n63447), .ZN(n25564) );
  INV_X1 U30035 ( .A(n25564), .ZN(p_wishbone_bd_ram_n25302) );
  INV_X1 U30036 ( .A(n63446), .ZN(n25566) );
  INV_X1 U30037 ( .A(n25566), .ZN(p_wishbone_bd_ram_n25301) );
  INV_X1 U30038 ( .A(n63445), .ZN(n25568) );
  INV_X1 U30039 ( .A(n25568), .ZN(p_wishbone_bd_ram_n25300) );
  INV_X1 U30040 ( .A(n63444), .ZN(n25570) );
  INV_X1 U30041 ( .A(n25570), .ZN(p_wishbone_bd_ram_n25299) );
  INV_X1 U30042 ( .A(n63443), .ZN(n25572) );
  INV_X1 U30043 ( .A(n25572), .ZN(p_wishbone_bd_ram_n25298) );
  INV_X1 U30044 ( .A(n63442), .ZN(n25574) );
  INV_X1 U30045 ( .A(n25574), .ZN(p_wishbone_bd_ram_n25297) );
  INV_X1 U30046 ( .A(n63441), .ZN(n25576) );
  INV_X1 U30047 ( .A(n25576), .ZN(p_wishbone_bd_ram_n25296) );
  INV_X1 U30048 ( .A(n63440), .ZN(n25578) );
  INV_X1 U30049 ( .A(n25578), .ZN(p_wishbone_bd_ram_n25295) );
  INV_X1 U30050 ( .A(n63439), .ZN(n25580) );
  INV_X1 U30051 ( .A(n25580), .ZN(p_wishbone_bd_ram_n25294) );
  INV_X1 U30052 ( .A(n63438), .ZN(n25582) );
  INV_X1 U30053 ( .A(n25582), .ZN(p_wishbone_bd_ram_n25293) );
  INV_X1 U30054 ( .A(n63437), .ZN(n25584) );
  INV_X1 U30055 ( .A(n25584), .ZN(p_wishbone_bd_ram_n25292) );
  INV_X1 U30056 ( .A(n63436), .ZN(n25586) );
  INV_X1 U30057 ( .A(n25586), .ZN(p_wishbone_bd_ram_n25291) );
  INV_X1 U30058 ( .A(n63435), .ZN(n25588) );
  INV_X1 U30059 ( .A(n25588), .ZN(p_wishbone_bd_ram_n25290) );
  INV_X1 U30060 ( .A(n63434), .ZN(n25590) );
  INV_X1 U30061 ( .A(n25590), .ZN(p_wishbone_bd_ram_n25289) );
  INV_X1 U30062 ( .A(n63433), .ZN(n25592) );
  INV_X1 U30063 ( .A(n25592), .ZN(p_wishbone_bd_ram_n25288) );
  INV_X1 U30064 ( .A(n63432), .ZN(n25594) );
  INV_X1 U30065 ( .A(n25594), .ZN(p_wishbone_bd_ram_n25287) );
  INV_X1 U30066 ( .A(n63431), .ZN(n25596) );
  INV_X1 U30067 ( .A(n25596), .ZN(p_wishbone_bd_ram_n25286) );
  INV_X1 U30068 ( .A(n63430), .ZN(n25598) );
  INV_X1 U30069 ( .A(n25598), .ZN(p_wishbone_bd_ram_n25285) );
  INV_X1 U30070 ( .A(n63429), .ZN(n25600) );
  INV_X1 U30071 ( .A(n25600), .ZN(p_wishbone_bd_ram_n25284) );
  INV_X1 U30072 ( .A(n63428), .ZN(n25602) );
  INV_X1 U30073 ( .A(n25602), .ZN(p_wishbone_bd_ram_n25283) );
  INV_X1 U30074 ( .A(n63427), .ZN(n25604) );
  INV_X1 U30075 ( .A(n25604), .ZN(p_wishbone_bd_ram_n25282) );
  INV_X1 U30076 ( .A(n63426), .ZN(n25606) );
  INV_X1 U30077 ( .A(n25606), .ZN(p_wishbone_bd_ram_n25281) );
  INV_X1 U30078 ( .A(n63425), .ZN(n25608) );
  INV_X1 U30079 ( .A(n25608), .ZN(p_wishbone_bd_ram_n25280) );
  INV_X1 U30080 ( .A(n63424), .ZN(n25610) );
  INV_X1 U30081 ( .A(n25610), .ZN(p_wishbone_bd_ram_n25279) );
  INV_X1 U30082 ( .A(n63423), .ZN(n25612) );
  INV_X1 U30083 ( .A(n25612), .ZN(p_wishbone_bd_ram_n25278) );
  INV_X1 U30084 ( .A(n63422), .ZN(n25614) );
  INV_X1 U30085 ( .A(n25614), .ZN(p_wishbone_bd_ram_n25277) );
  INV_X1 U30086 ( .A(n63421), .ZN(n25616) );
  INV_X1 U30087 ( .A(n25616), .ZN(p_wishbone_bd_ram_n25276) );
  INV_X1 U30088 ( .A(n63420), .ZN(n25618) );
  INV_X1 U30089 ( .A(n25618), .ZN(p_wishbone_bd_ram_n25275) );
  INV_X1 U30090 ( .A(n63419), .ZN(n25620) );
  INV_X1 U30091 ( .A(n25620), .ZN(p_wishbone_bd_ram_n25274) );
  INV_X1 U30092 ( .A(n63418), .ZN(n25622) );
  INV_X1 U30093 ( .A(n25622), .ZN(p_wishbone_bd_ram_n25273) );
  INV_X1 U30094 ( .A(n63417), .ZN(n25624) );
  INV_X1 U30095 ( .A(n25624), .ZN(p_wishbone_bd_ram_n25272) );
  INV_X1 U30096 ( .A(n63416), .ZN(n25626) );
  INV_X1 U30097 ( .A(n25626), .ZN(p_wishbone_bd_ram_n25271) );
  INV_X1 U30098 ( .A(n63415), .ZN(n25628) );
  INV_X1 U30099 ( .A(n25628), .ZN(p_wishbone_bd_ram_n25270) );
  INV_X1 U30100 ( .A(n63414), .ZN(n25630) );
  INV_X1 U30101 ( .A(n25630), .ZN(p_wishbone_bd_ram_n25269) );
  INV_X1 U30102 ( .A(n63413), .ZN(n25632) );
  INV_X1 U30103 ( .A(n25632), .ZN(p_wishbone_bd_ram_n25268) );
  INV_X1 U30104 ( .A(n63412), .ZN(n25634) );
  INV_X1 U30105 ( .A(n25634), .ZN(p_wishbone_bd_ram_n25267) );
  INV_X1 U30106 ( .A(n63411), .ZN(n25636) );
  INV_X1 U30107 ( .A(n25636), .ZN(p_wishbone_bd_ram_n25266) );
  INV_X1 U30108 ( .A(n63410), .ZN(n25638) );
  INV_X1 U30109 ( .A(n25638), .ZN(p_wishbone_bd_ram_n25265) );
  INV_X1 U30110 ( .A(n63409), .ZN(n25640) );
  INV_X1 U30111 ( .A(n25640), .ZN(p_wishbone_bd_ram_n25263) );
  INV_X1 U30112 ( .A(n63408), .ZN(n25642) );
  INV_X1 U30113 ( .A(n25642), .ZN(p_wishbone_bd_ram_n25261) );
  INV_X1 U30114 ( .A(n63407), .ZN(n25644) );
  INV_X1 U30115 ( .A(n25644), .ZN(p_wishbone_bd_ram_n25260) );
  INV_X1 U30116 ( .A(n63406), .ZN(n25646) );
  INV_X1 U30117 ( .A(n25646), .ZN(p_wishbone_bd_ram_n25258) );
  INV_X1 U30118 ( .A(n63405), .ZN(n25648) );
  INV_X1 U30119 ( .A(n25648), .ZN(p_wishbone_bd_ram_n25256) );
  INV_X1 U30120 ( .A(n63404), .ZN(n25650) );
  INV_X1 U30121 ( .A(n25650), .ZN(p_wishbone_bd_ram_n25255) );
  INV_X1 U30122 ( .A(n63403), .ZN(n25652) );
  INV_X1 U30123 ( .A(n25652), .ZN(p_wishbone_bd_ram_n25254) );
  INV_X1 U30124 ( .A(n63402), .ZN(n25654) );
  INV_X1 U30125 ( .A(n25654), .ZN(p_wishbone_bd_ram_n25253) );
  INV_X1 U30126 ( .A(n63401), .ZN(n25656) );
  INV_X1 U30127 ( .A(n25656), .ZN(p_wishbone_bd_ram_n25252) );
  INV_X1 U30128 ( .A(n63400), .ZN(n25658) );
  INV_X1 U30129 ( .A(n25658), .ZN(p_wishbone_bd_ram_n25251) );
  INV_X1 U30130 ( .A(n63399), .ZN(n25660) );
  INV_X1 U30131 ( .A(n25660), .ZN(p_wishbone_bd_ram_n25250) );
  INV_X1 U30132 ( .A(n63398), .ZN(n25662) );
  INV_X1 U30133 ( .A(n25662), .ZN(p_wishbone_bd_ram_n25249) );
  INV_X1 U30134 ( .A(n63397), .ZN(n25664) );
  INV_X1 U30135 ( .A(n25664), .ZN(p_wishbone_bd_ram_n25248) );
  INV_X1 U30136 ( .A(n63396), .ZN(n25666) );
  INV_X1 U30137 ( .A(n25666), .ZN(p_wishbone_bd_ram_n25247) );
  INV_X1 U30138 ( .A(n63395), .ZN(n25668) );
  INV_X1 U30139 ( .A(n25668), .ZN(p_wishbone_bd_ram_n25246) );
  INV_X1 U30140 ( .A(n63394), .ZN(n25670) );
  INV_X1 U30141 ( .A(n25670), .ZN(p_wishbone_bd_ram_n25245) );
  INV_X1 U30142 ( .A(n63393), .ZN(n25672) );
  INV_X1 U30143 ( .A(n25672), .ZN(p_wishbone_bd_ram_n25244) );
  INV_X1 U30144 ( .A(n63392), .ZN(n25674) );
  INV_X1 U30145 ( .A(n25674), .ZN(p_wishbone_bd_ram_n25243) );
  INV_X1 U30146 ( .A(n63391), .ZN(n25676) );
  INV_X1 U30147 ( .A(n25676), .ZN(p_wishbone_bd_ram_n25242) );
  INV_X1 U30148 ( .A(n63390), .ZN(n25678) );
  INV_X1 U30149 ( .A(n25678), .ZN(p_wishbone_bd_ram_n25241) );
  INV_X1 U30150 ( .A(n63389), .ZN(n25680) );
  INV_X1 U30151 ( .A(n25680), .ZN(p_wishbone_bd_ram_n25240) );
  INV_X1 U30152 ( .A(n63388), .ZN(n25682) );
  INV_X1 U30153 ( .A(n25682), .ZN(p_wishbone_bd_ram_n25239) );
  INV_X1 U30154 ( .A(n63387), .ZN(n25684) );
  INV_X1 U30155 ( .A(n25684), .ZN(p_wishbone_bd_ram_n25238) );
  INV_X1 U30156 ( .A(n63386), .ZN(n25686) );
  INV_X1 U30157 ( .A(n25686), .ZN(p_wishbone_bd_ram_n25237) );
  INV_X1 U30158 ( .A(n63385), .ZN(n25688) );
  INV_X1 U30159 ( .A(n25688), .ZN(p_wishbone_bd_ram_n25236) );
  INV_X1 U30160 ( .A(n63384), .ZN(n25690) );
  INV_X1 U30161 ( .A(n25690), .ZN(p_wishbone_bd_ram_n25235) );
  INV_X1 U30162 ( .A(n63383), .ZN(n25692) );
  INV_X1 U30163 ( .A(n25692), .ZN(p_wishbone_bd_ram_n25234) );
  INV_X1 U30164 ( .A(n63382), .ZN(n25694) );
  INV_X1 U30165 ( .A(n25694), .ZN(p_wishbone_bd_ram_n25233) );
  INV_X1 U30166 ( .A(n63381), .ZN(n25696) );
  INV_X1 U30167 ( .A(n25696), .ZN(p_wishbone_bd_ram_n25232) );
  INV_X1 U30168 ( .A(n63380), .ZN(n25698) );
  INV_X1 U30169 ( .A(n25698), .ZN(p_wishbone_bd_ram_n25231) );
  INV_X1 U30170 ( .A(n63379), .ZN(n25700) );
  INV_X1 U30171 ( .A(n25700), .ZN(p_wishbone_bd_ram_n25230) );
  INV_X1 U30172 ( .A(n63378), .ZN(n25702) );
  INV_X1 U30173 ( .A(n25702), .ZN(p_wishbone_bd_ram_n25229) );
  INV_X1 U30174 ( .A(n63377), .ZN(n25704) );
  INV_X1 U30175 ( .A(n25704), .ZN(p_wishbone_bd_ram_n25228) );
  INV_X1 U30176 ( .A(n63376), .ZN(n25706) );
  INV_X1 U30177 ( .A(n25706), .ZN(p_wishbone_bd_ram_n25227) );
  INV_X1 U30178 ( .A(n63375), .ZN(n25708) );
  INV_X1 U30179 ( .A(n25708), .ZN(p_wishbone_bd_ram_n25226) );
  INV_X1 U30180 ( .A(n63374), .ZN(n25710) );
  INV_X1 U30181 ( .A(n25710), .ZN(p_wishbone_bd_ram_n25225) );
  INV_X1 U30182 ( .A(n63373), .ZN(n25712) );
  INV_X1 U30183 ( .A(n25712), .ZN(p_wishbone_bd_ram_n25224) );
  INV_X1 U30184 ( .A(n63372), .ZN(n25714) );
  INV_X1 U30185 ( .A(n25714), .ZN(p_wishbone_bd_ram_n25223) );
  INV_X1 U30186 ( .A(n63371), .ZN(n25716) );
  INV_X1 U30187 ( .A(n25716), .ZN(p_wishbone_bd_ram_n25222) );
  INV_X1 U30188 ( .A(n63370), .ZN(n25718) );
  INV_X1 U30189 ( .A(n25718), .ZN(p_wishbone_bd_ram_n25221) );
  INV_X1 U30190 ( .A(n63369), .ZN(n25720) );
  INV_X1 U30191 ( .A(n25720), .ZN(p_wishbone_bd_ram_n25220) );
  INV_X1 U30192 ( .A(n63368), .ZN(n25722) );
  INV_X1 U30193 ( .A(n25722), .ZN(p_wishbone_bd_ram_n25219) );
  INV_X1 U30194 ( .A(n63367), .ZN(n25724) );
  INV_X1 U30195 ( .A(n25724), .ZN(p_wishbone_bd_ram_n25218) );
  INV_X1 U30196 ( .A(n63366), .ZN(n25726) );
  INV_X1 U30197 ( .A(n25726), .ZN(p_wishbone_bd_ram_n25217) );
  INV_X1 U30198 ( .A(n63365), .ZN(n25728) );
  INV_X1 U30199 ( .A(n25728), .ZN(p_wishbone_bd_ram_n25216) );
  INV_X1 U30200 ( .A(n63364), .ZN(n25730) );
  INV_X1 U30201 ( .A(n25730), .ZN(p_wishbone_bd_ram_n25215) );
  INV_X1 U30202 ( .A(n63363), .ZN(n25732) );
  INV_X1 U30203 ( .A(n25732), .ZN(p_wishbone_bd_ram_n25214) );
  INV_X1 U30204 ( .A(n63362), .ZN(n25734) );
  INV_X1 U30205 ( .A(n25734), .ZN(p_wishbone_bd_ram_n25213) );
  INV_X1 U30206 ( .A(n63361), .ZN(n25736) );
  INV_X1 U30207 ( .A(n25736), .ZN(p_wishbone_bd_ram_n25212) );
  INV_X1 U30208 ( .A(n63360), .ZN(n25738) );
  INV_X1 U30209 ( .A(n25738), .ZN(p_wishbone_bd_ram_n25211) );
  INV_X1 U30210 ( .A(n63359), .ZN(n25740) );
  INV_X1 U30211 ( .A(n25740), .ZN(p_wishbone_bd_ram_n25210) );
  INV_X1 U30212 ( .A(n63358), .ZN(n25742) );
  INV_X1 U30213 ( .A(n25742), .ZN(p_wishbone_bd_ram_n25209) );
  INV_X1 U30214 ( .A(n63357), .ZN(n25744) );
  INV_X1 U30215 ( .A(n25744), .ZN(p_wishbone_bd_ram_n25207) );
  INV_X1 U30216 ( .A(n63356), .ZN(n25746) );
  INV_X1 U30217 ( .A(n25746), .ZN(p_wishbone_bd_ram_n25205) );
  INV_X1 U30218 ( .A(n63355), .ZN(n25748) );
  INV_X1 U30219 ( .A(n25748), .ZN(p_wishbone_bd_ram_n25204) );
  INV_X1 U30220 ( .A(n63354), .ZN(n25750) );
  INV_X1 U30221 ( .A(n25750), .ZN(p_wishbone_bd_ram_n25202) );
  INV_X1 U30222 ( .A(n63353), .ZN(n25752) );
  INV_X1 U30223 ( .A(n25752), .ZN(p_wishbone_bd_ram_n25200) );
  INV_X1 U30224 ( .A(n63352), .ZN(n25754) );
  INV_X1 U30225 ( .A(n25754), .ZN(p_wishbone_bd_ram_n25199) );
  INV_X1 U30226 ( .A(n63351), .ZN(n25756) );
  INV_X1 U30227 ( .A(n25756), .ZN(p_wishbone_bd_ram_n25198) );
  INV_X1 U30228 ( .A(n63350), .ZN(n25758) );
  INV_X1 U30229 ( .A(n25758), .ZN(p_wishbone_bd_ram_n25197) );
  INV_X1 U30230 ( .A(n63349), .ZN(n25760) );
  INV_X1 U30231 ( .A(n25760), .ZN(p_wishbone_bd_ram_n25196) );
  INV_X1 U30232 ( .A(n63348), .ZN(n25762) );
  INV_X1 U30233 ( .A(n25762), .ZN(p_wishbone_bd_ram_n25195) );
  INV_X1 U30234 ( .A(n63347), .ZN(n25764) );
  INV_X1 U30235 ( .A(n25764), .ZN(p_wishbone_bd_ram_n25194) );
  INV_X1 U30236 ( .A(n63346), .ZN(n25766) );
  INV_X1 U30237 ( .A(n25766), .ZN(p_wishbone_bd_ram_n25193) );
  INV_X1 U30238 ( .A(n63345), .ZN(n25768) );
  INV_X1 U30239 ( .A(n25768), .ZN(p_wishbone_bd_ram_n25192) );
  INV_X1 U30240 ( .A(n63344), .ZN(n25770) );
  INV_X1 U30241 ( .A(n25770), .ZN(p_wishbone_bd_ram_n25191) );
  INV_X1 U30242 ( .A(n63343), .ZN(n25772) );
  INV_X1 U30243 ( .A(n25772), .ZN(p_wishbone_bd_ram_n25190) );
  INV_X1 U30244 ( .A(n63342), .ZN(n25774) );
  INV_X1 U30245 ( .A(n25774), .ZN(p_wishbone_bd_ram_n25189) );
  INV_X1 U30246 ( .A(n63341), .ZN(n25776) );
  INV_X1 U30247 ( .A(n25776), .ZN(p_wishbone_bd_ram_n25188) );
  INV_X1 U30248 ( .A(n63340), .ZN(n25778) );
  INV_X1 U30249 ( .A(n25778), .ZN(p_wishbone_bd_ram_n25187) );
  INV_X1 U30250 ( .A(n63339), .ZN(n25780) );
  INV_X1 U30251 ( .A(n25780), .ZN(p_wishbone_bd_ram_n25186) );
  INV_X1 U30252 ( .A(n63338), .ZN(n25782) );
  INV_X1 U30253 ( .A(n25782), .ZN(p_wishbone_bd_ram_n25185) );
  INV_X1 U30254 ( .A(n63337), .ZN(n25784) );
  INV_X1 U30255 ( .A(n25784), .ZN(p_wishbone_bd_ram_n25184) );
  INV_X1 U30256 ( .A(n63336), .ZN(n25786) );
  INV_X1 U30257 ( .A(n25786), .ZN(p_wishbone_bd_ram_n25183) );
  INV_X1 U30258 ( .A(n63335), .ZN(n25788) );
  INV_X1 U30259 ( .A(n25788), .ZN(p_wishbone_bd_ram_n25182) );
  INV_X1 U30260 ( .A(n63334), .ZN(n25790) );
  INV_X1 U30261 ( .A(n25790), .ZN(p_wishbone_bd_ram_n25181) );
  INV_X1 U30262 ( .A(n63333), .ZN(n25792) );
  INV_X1 U30263 ( .A(n25792), .ZN(p_wishbone_bd_ram_n25180) );
  INV_X1 U30264 ( .A(n63332), .ZN(n25794) );
  INV_X1 U30265 ( .A(n25794), .ZN(p_wishbone_bd_ram_n25179) );
  INV_X1 U30266 ( .A(n63331), .ZN(n25796) );
  INV_X1 U30267 ( .A(n25796), .ZN(p_wishbone_bd_ram_n25178) );
  INV_X1 U30268 ( .A(n63330), .ZN(n25798) );
  INV_X1 U30269 ( .A(n25798), .ZN(p_wishbone_bd_ram_n25177) );
  INV_X1 U30270 ( .A(n63329), .ZN(n25800) );
  INV_X1 U30271 ( .A(n25800), .ZN(p_wishbone_bd_ram_n25176) );
  INV_X1 U30272 ( .A(n63328), .ZN(n25802) );
  INV_X1 U30273 ( .A(n25802), .ZN(p_wishbone_bd_ram_n25175) );
  INV_X1 U30274 ( .A(n63327), .ZN(n25804) );
  INV_X1 U30275 ( .A(n25804), .ZN(p_wishbone_bd_ram_n25174) );
  INV_X1 U30276 ( .A(n63326), .ZN(n25806) );
  INV_X1 U30277 ( .A(n25806), .ZN(p_wishbone_bd_ram_n25173) );
  INV_X1 U30278 ( .A(n63325), .ZN(n25808) );
  INV_X1 U30279 ( .A(n25808), .ZN(p_wishbone_bd_ram_n25172) );
  INV_X1 U30280 ( .A(n63324), .ZN(n25810) );
  INV_X1 U30281 ( .A(n25810), .ZN(p_wishbone_bd_ram_n25171) );
  INV_X1 U30282 ( .A(n63323), .ZN(n25812) );
  INV_X1 U30283 ( .A(n25812), .ZN(p_wishbone_bd_ram_n25170) );
  INV_X1 U30284 ( .A(n63322), .ZN(n25814) );
  INV_X1 U30285 ( .A(n25814), .ZN(p_wishbone_bd_ram_n25169) );
  INV_X1 U30286 ( .A(n63321), .ZN(n25816) );
  INV_X1 U30287 ( .A(n25816), .ZN(p_wishbone_bd_ram_n25168) );
  INV_X1 U30288 ( .A(n63320), .ZN(n25818) );
  INV_X1 U30289 ( .A(n25818), .ZN(p_wishbone_bd_ram_n25167) );
  INV_X1 U30290 ( .A(n63319), .ZN(n25820) );
  INV_X1 U30291 ( .A(n25820), .ZN(p_wishbone_bd_ram_n25166) );
  INV_X1 U30292 ( .A(n63318), .ZN(n25822) );
  INV_X1 U30293 ( .A(n25822), .ZN(p_wishbone_bd_ram_n25165) );
  INV_X1 U30294 ( .A(n63317), .ZN(n25824) );
  INV_X1 U30295 ( .A(n25824), .ZN(p_wishbone_bd_ram_n25164) );
  INV_X1 U30296 ( .A(n63316), .ZN(n25826) );
  INV_X1 U30297 ( .A(n25826), .ZN(p_wishbone_bd_ram_n25163) );
  INV_X1 U30298 ( .A(n63315), .ZN(n25828) );
  INV_X1 U30299 ( .A(n25828), .ZN(p_wishbone_bd_ram_n25162) );
  INV_X1 U30300 ( .A(n63314), .ZN(n25830) );
  INV_X1 U30301 ( .A(n25830), .ZN(p_wishbone_bd_ram_n25161) );
  INV_X1 U30302 ( .A(n63313), .ZN(n25832) );
  INV_X1 U30303 ( .A(n25832), .ZN(p_wishbone_bd_ram_n25160) );
  INV_X1 U30304 ( .A(n63312), .ZN(n25834) );
  INV_X1 U30305 ( .A(n25834), .ZN(p_wishbone_bd_ram_n25159) );
  INV_X1 U30306 ( .A(n63311), .ZN(n25836) );
  INV_X1 U30307 ( .A(n25836), .ZN(p_wishbone_bd_ram_n25158) );
  INV_X1 U30308 ( .A(n63310), .ZN(n25838) );
  INV_X1 U30309 ( .A(n25838), .ZN(p_wishbone_bd_ram_n25157) );
  INV_X1 U30310 ( .A(n63309), .ZN(n25840) );
  INV_X1 U30311 ( .A(n25840), .ZN(p_wishbone_bd_ram_n25156) );
  INV_X1 U30312 ( .A(n63308), .ZN(n25842) );
  INV_X1 U30313 ( .A(n25842), .ZN(p_wishbone_bd_ram_n25155) );
  INV_X1 U30314 ( .A(n63307), .ZN(n25844) );
  INV_X1 U30315 ( .A(n25844), .ZN(p_wishbone_bd_ram_n25154) );
  INV_X1 U30316 ( .A(n63306), .ZN(n25846) );
  INV_X1 U30317 ( .A(n25846), .ZN(p_wishbone_bd_ram_n25153) );
  INV_X1 U30318 ( .A(n63305), .ZN(n25848) );
  INV_X1 U30319 ( .A(n25848), .ZN(p_wishbone_bd_ram_n25152) );
  INV_X1 U30320 ( .A(n63304), .ZN(n25850) );
  INV_X1 U30321 ( .A(n25850), .ZN(p_wishbone_bd_ram_n25151) );
  INV_X1 U30322 ( .A(n63303), .ZN(n25852) );
  INV_X1 U30323 ( .A(n25852), .ZN(p_wishbone_bd_ram_n25150) );
  INV_X1 U30324 ( .A(n63302), .ZN(n25854) );
  INV_X1 U30325 ( .A(n25854), .ZN(p_wishbone_bd_ram_n25149) );
  INV_X1 U30326 ( .A(n63301), .ZN(n25856) );
  INV_X1 U30327 ( .A(n25856), .ZN(p_wishbone_bd_ram_n25148) );
  INV_X1 U30328 ( .A(n63300), .ZN(n25858) );
  INV_X1 U30329 ( .A(n25858), .ZN(p_wishbone_bd_ram_n25147) );
  INV_X1 U30330 ( .A(n63299), .ZN(n25860) );
  INV_X1 U30331 ( .A(n25860), .ZN(p_wishbone_bd_ram_n25146) );
  INV_X1 U30332 ( .A(n63298), .ZN(n25862) );
  INV_X1 U30333 ( .A(n25862), .ZN(p_wishbone_bd_ram_n25145) );
  INV_X1 U30334 ( .A(n63297), .ZN(n25864) );
  INV_X1 U30335 ( .A(n25864), .ZN(p_wishbone_bd_ram_n25144) );
  INV_X1 U30336 ( .A(n63296), .ZN(n25866) );
  INV_X1 U30337 ( .A(n25866), .ZN(p_wishbone_bd_ram_n25143) );
  INV_X1 U30338 ( .A(n63295), .ZN(n25868) );
  INV_X1 U30339 ( .A(n25868), .ZN(p_wishbone_bd_ram_n25142) );
  INV_X1 U30340 ( .A(n63294), .ZN(n25870) );
  INV_X1 U30341 ( .A(n25870), .ZN(p_wishbone_bd_ram_n25141) );
  INV_X1 U30342 ( .A(n63293), .ZN(n25872) );
  INV_X1 U30343 ( .A(n25872), .ZN(p_wishbone_bd_ram_n25140) );
  INV_X1 U30344 ( .A(n63292), .ZN(n25874) );
  INV_X1 U30345 ( .A(n25874), .ZN(p_wishbone_bd_ram_n25139) );
  INV_X1 U30346 ( .A(n63291), .ZN(n25876) );
  INV_X1 U30347 ( .A(n25876), .ZN(p_wishbone_bd_ram_n25138) );
  INV_X1 U30348 ( .A(n63290), .ZN(n25878) );
  INV_X1 U30349 ( .A(n25878), .ZN(p_wishbone_bd_ram_n25137) );
  INV_X1 U30350 ( .A(n63289), .ZN(n25880) );
  INV_X1 U30351 ( .A(n25880), .ZN(p_wishbone_bd_ram_n25135) );
  INV_X1 U30352 ( .A(n63288), .ZN(n25882) );
  INV_X1 U30353 ( .A(n25882), .ZN(p_wishbone_bd_ram_n25133) );
  INV_X1 U30354 ( .A(n63287), .ZN(n25884) );
  INV_X1 U30355 ( .A(n25884), .ZN(p_wishbone_bd_ram_n25132) );
  INV_X1 U30356 ( .A(n63286), .ZN(n25886) );
  INV_X1 U30357 ( .A(n25886), .ZN(p_wishbone_bd_ram_n25130) );
  INV_X1 U30358 ( .A(n63285), .ZN(n25888) );
  INV_X1 U30359 ( .A(n25888), .ZN(p_wishbone_bd_ram_n25128) );
  INV_X1 U30360 ( .A(n63284), .ZN(n25890) );
  INV_X1 U30361 ( .A(n25890), .ZN(p_wishbone_bd_ram_n25127) );
  INV_X1 U30362 ( .A(n63283), .ZN(n25892) );
  INV_X1 U30363 ( .A(n25892), .ZN(p_wishbone_bd_ram_n25126) );
  INV_X1 U30364 ( .A(n63282), .ZN(n25894) );
  INV_X1 U30365 ( .A(n25894), .ZN(p_wishbone_bd_ram_n25125) );
  INV_X1 U30366 ( .A(n63281), .ZN(n25896) );
  INV_X1 U30367 ( .A(n25896), .ZN(p_wishbone_bd_ram_n25124) );
  INV_X1 U30368 ( .A(n63280), .ZN(n25898) );
  INV_X1 U30369 ( .A(n25898), .ZN(p_wishbone_bd_ram_n25123) );
  INV_X1 U30370 ( .A(n63279), .ZN(n25900) );
  INV_X1 U30371 ( .A(n25900), .ZN(p_wishbone_bd_ram_n25122) );
  INV_X1 U30372 ( .A(n63278), .ZN(n25902) );
  INV_X1 U30373 ( .A(n25902), .ZN(p_wishbone_bd_ram_n25121) );
  INV_X1 U30374 ( .A(n63277), .ZN(n25904) );
  INV_X1 U30375 ( .A(n25904), .ZN(p_wishbone_bd_ram_n25120) );
  INV_X1 U30376 ( .A(n63276), .ZN(n25906) );
  INV_X1 U30377 ( .A(n25906), .ZN(p_wishbone_bd_ram_n25119) );
  INV_X1 U30378 ( .A(n63275), .ZN(n25908) );
  INV_X1 U30379 ( .A(n25908), .ZN(p_wishbone_bd_ram_n25118) );
  INV_X1 U30380 ( .A(n63274), .ZN(n25910) );
  INV_X1 U30381 ( .A(n25910), .ZN(p_wishbone_bd_ram_n25117) );
  INV_X1 U30382 ( .A(n63273), .ZN(n25912) );
  INV_X1 U30383 ( .A(n25912), .ZN(p_wishbone_bd_ram_n25116) );
  INV_X1 U30384 ( .A(n63272), .ZN(n25914) );
  INV_X1 U30385 ( .A(n25914), .ZN(p_wishbone_bd_ram_n25115) );
  INV_X1 U30386 ( .A(n63271), .ZN(n25916) );
  INV_X1 U30387 ( .A(n25916), .ZN(p_wishbone_bd_ram_n25114) );
  INV_X1 U30388 ( .A(n63270), .ZN(n25918) );
  INV_X1 U30389 ( .A(n25918), .ZN(p_wishbone_bd_ram_n25113) );
  INV_X1 U30390 ( .A(n63269), .ZN(n25920) );
  INV_X1 U30391 ( .A(n25920), .ZN(p_wishbone_bd_ram_n25112) );
  INV_X1 U30392 ( .A(n63268), .ZN(n25922) );
  INV_X1 U30393 ( .A(n25922), .ZN(p_wishbone_bd_ram_n25111) );
  INV_X1 U30394 ( .A(n63267), .ZN(n25924) );
  INV_X1 U30395 ( .A(n25924), .ZN(p_wishbone_bd_ram_n25110) );
  INV_X1 U30396 ( .A(n63266), .ZN(n25926) );
  INV_X1 U30397 ( .A(n25926), .ZN(p_wishbone_bd_ram_n25109) );
  INV_X1 U30398 ( .A(n63265), .ZN(n25928) );
  INV_X1 U30399 ( .A(n25928), .ZN(p_wishbone_bd_ram_n25108) );
  INV_X1 U30400 ( .A(n63264), .ZN(n25930) );
  INV_X1 U30401 ( .A(n25930), .ZN(p_wishbone_bd_ram_n25107) );
  INV_X1 U30402 ( .A(n63263), .ZN(n25932) );
  INV_X1 U30403 ( .A(n25932), .ZN(p_wishbone_bd_ram_n25106) );
  INV_X1 U30404 ( .A(n63262), .ZN(n25934) );
  INV_X1 U30405 ( .A(n25934), .ZN(p_wishbone_bd_ram_n25105) );
  INV_X1 U30406 ( .A(n63261), .ZN(n25936) );
  INV_X1 U30407 ( .A(n25936), .ZN(p_wishbone_bd_ram_n25104) );
  INV_X1 U30408 ( .A(n63260), .ZN(n25938) );
  INV_X1 U30409 ( .A(n25938), .ZN(p_wishbone_bd_ram_n25103) );
  INV_X1 U30410 ( .A(n63259), .ZN(n25940) );
  INV_X1 U30411 ( .A(n25940), .ZN(p_wishbone_bd_ram_n25102) );
  INV_X1 U30412 ( .A(n63258), .ZN(n25942) );
  INV_X1 U30413 ( .A(n25942), .ZN(p_wishbone_bd_ram_n25101) );
  INV_X1 U30414 ( .A(n63257), .ZN(n25944) );
  INV_X1 U30415 ( .A(n25944), .ZN(p_wishbone_bd_ram_n25100) );
  INV_X1 U30416 ( .A(n63256), .ZN(n25946) );
  INV_X1 U30417 ( .A(n25946), .ZN(p_wishbone_bd_ram_n25099) );
  INV_X1 U30418 ( .A(n63255), .ZN(n25948) );
  INV_X1 U30419 ( .A(n25948), .ZN(p_wishbone_bd_ram_n25098) );
  INV_X1 U30420 ( .A(n63254), .ZN(n25950) );
  INV_X1 U30421 ( .A(n25950), .ZN(p_wishbone_bd_ram_n25097) );
  INV_X1 U30422 ( .A(n63253), .ZN(n25952) );
  INV_X1 U30423 ( .A(n25952), .ZN(p_wishbone_bd_ram_n25096) );
  INV_X1 U30424 ( .A(n63252), .ZN(n25954) );
  INV_X1 U30425 ( .A(n25954), .ZN(p_wishbone_bd_ram_n25095) );
  INV_X1 U30426 ( .A(n63251), .ZN(n25956) );
  INV_X1 U30427 ( .A(n25956), .ZN(p_wishbone_bd_ram_n25094) );
  INV_X1 U30428 ( .A(n63250), .ZN(n25958) );
  INV_X1 U30429 ( .A(n25958), .ZN(p_wishbone_bd_ram_n25093) );
  INV_X1 U30430 ( .A(n63249), .ZN(n25960) );
  INV_X1 U30431 ( .A(n25960), .ZN(p_wishbone_bd_ram_n25092) );
  INV_X1 U30432 ( .A(n63248), .ZN(n25962) );
  INV_X1 U30433 ( .A(n25962), .ZN(p_wishbone_bd_ram_n25091) );
  INV_X1 U30434 ( .A(n63247), .ZN(n25964) );
  INV_X1 U30435 ( .A(n25964), .ZN(p_wishbone_bd_ram_n25090) );
  INV_X1 U30436 ( .A(n63246), .ZN(n25966) );
  INV_X1 U30437 ( .A(n25966), .ZN(p_wishbone_bd_ram_n25089) );
  INV_X1 U30438 ( .A(n63245), .ZN(n25968) );
  INV_X1 U30439 ( .A(n25968), .ZN(p_wishbone_bd_ram_n25088) );
  INV_X1 U30440 ( .A(n63244), .ZN(n25970) );
  INV_X1 U30441 ( .A(n25970), .ZN(p_wishbone_bd_ram_n25087) );
  INV_X1 U30442 ( .A(n63243), .ZN(n25972) );
  INV_X1 U30443 ( .A(n25972), .ZN(p_wishbone_bd_ram_n25086) );
  INV_X1 U30444 ( .A(n63242), .ZN(n25974) );
  INV_X1 U30445 ( .A(n25974), .ZN(p_wishbone_bd_ram_n25085) );
  INV_X1 U30446 ( .A(n63241), .ZN(n25976) );
  INV_X1 U30447 ( .A(n25976), .ZN(p_wishbone_bd_ram_n25084) );
  INV_X1 U30448 ( .A(n63240), .ZN(n25978) );
  INV_X1 U30449 ( .A(n25978), .ZN(p_wishbone_bd_ram_n25083) );
  INV_X1 U30450 ( .A(n63239), .ZN(n25980) );
  INV_X1 U30451 ( .A(n25980), .ZN(p_wishbone_bd_ram_n25082) );
  INV_X1 U30452 ( .A(n63238), .ZN(n25982) );
  INV_X1 U30453 ( .A(n25982), .ZN(p_wishbone_bd_ram_n25081) );
  INV_X1 U30454 ( .A(n63237), .ZN(n25984) );
  INV_X1 U30455 ( .A(n25984), .ZN(p_wishbone_bd_ram_n25080) );
  INV_X1 U30456 ( .A(n63236), .ZN(n25986) );
  INV_X1 U30457 ( .A(n25986), .ZN(p_wishbone_bd_ram_n25079) );
  INV_X1 U30458 ( .A(n63235), .ZN(n25988) );
  INV_X1 U30459 ( .A(n25988), .ZN(p_wishbone_bd_ram_n25078) );
  INV_X1 U30460 ( .A(n63234), .ZN(n25990) );
  INV_X1 U30461 ( .A(n25990), .ZN(p_wishbone_bd_ram_n25077) );
  INV_X1 U30462 ( .A(n63233), .ZN(n25992) );
  INV_X1 U30463 ( .A(n25992), .ZN(p_wishbone_bd_ram_n25076) );
  INV_X1 U30464 ( .A(n63232), .ZN(n25994) );
  INV_X1 U30465 ( .A(n25994), .ZN(p_wishbone_bd_ram_n25075) );
  INV_X1 U30466 ( .A(n63231), .ZN(n25996) );
  INV_X1 U30467 ( .A(n25996), .ZN(p_wishbone_bd_ram_n25074) );
  INV_X1 U30468 ( .A(n63230), .ZN(n25998) );
  INV_X1 U30469 ( .A(n25998), .ZN(p_wishbone_bd_ram_n25073) );
  INV_X1 U30470 ( .A(n63229), .ZN(n26000) );
  INV_X1 U30471 ( .A(n26000), .ZN(p_wishbone_bd_ram_n25072) );
  INV_X1 U30472 ( .A(n63228), .ZN(n26002) );
  INV_X1 U30473 ( .A(n26002), .ZN(p_wishbone_bd_ram_n25071) );
  INV_X1 U30474 ( .A(n63227), .ZN(n26004) );
  INV_X1 U30475 ( .A(n26004), .ZN(p_wishbone_bd_ram_n25070) );
  INV_X1 U30476 ( .A(n63226), .ZN(n26006) );
  INV_X1 U30477 ( .A(n26006), .ZN(p_wishbone_bd_ram_n25069) );
  INV_X1 U30478 ( .A(n63225), .ZN(n26008) );
  INV_X1 U30479 ( .A(n26008), .ZN(p_wishbone_bd_ram_n25068) );
  INV_X1 U30480 ( .A(n63224), .ZN(n26010) );
  INV_X1 U30481 ( .A(n26010), .ZN(p_wishbone_bd_ram_n25067) );
  INV_X1 U30482 ( .A(n63223), .ZN(n26012) );
  INV_X1 U30483 ( .A(n26012), .ZN(p_wishbone_bd_ram_n25066) );
  INV_X1 U30484 ( .A(n63222), .ZN(n26014) );
  INV_X1 U30485 ( .A(n26014), .ZN(p_wishbone_bd_ram_n25065) );
  INV_X1 U30486 ( .A(n63221), .ZN(n26016) );
  INV_X1 U30487 ( .A(n26016), .ZN(p_wishbone_bd_ram_n25064) );
  INV_X1 U30488 ( .A(n63220), .ZN(n26018) );
  INV_X1 U30489 ( .A(n26018), .ZN(p_wishbone_bd_ram_n25063) );
  INV_X1 U30490 ( .A(n63219), .ZN(n26020) );
  INV_X1 U30491 ( .A(n26020), .ZN(p_wishbone_bd_ram_n25062) );
  INV_X1 U30492 ( .A(n63218), .ZN(n26022) );
  INV_X1 U30493 ( .A(n26022), .ZN(p_wishbone_bd_ram_n25061) );
  INV_X1 U30494 ( .A(n63217), .ZN(n26024) );
  INV_X1 U30495 ( .A(n26024), .ZN(p_wishbone_bd_ram_n25060) );
  INV_X1 U30496 ( .A(n63216), .ZN(n26026) );
  INV_X1 U30497 ( .A(n26026), .ZN(p_wishbone_bd_ram_n25059) );
  INV_X1 U30498 ( .A(n63215), .ZN(n26028) );
  INV_X1 U30499 ( .A(n26028), .ZN(p_wishbone_bd_ram_n25058) );
  INV_X1 U30500 ( .A(n63214), .ZN(n26030) );
  INV_X1 U30501 ( .A(n26030), .ZN(p_wishbone_bd_ram_n25057) );
  INV_X1 U30502 ( .A(n63213), .ZN(n26032) );
  INV_X1 U30503 ( .A(n26032), .ZN(p_wishbone_bd_ram_n25056) );
  INV_X1 U30504 ( .A(n63212), .ZN(n26034) );
  INV_X1 U30505 ( .A(n26034), .ZN(p_wishbone_bd_ram_n25055) );
  INV_X1 U30506 ( .A(n63211), .ZN(n26036) );
  INV_X1 U30507 ( .A(n26036), .ZN(p_wishbone_bd_ram_n25054) );
  INV_X1 U30508 ( .A(n63210), .ZN(n26038) );
  INV_X1 U30509 ( .A(n26038), .ZN(p_wishbone_bd_ram_n25053) );
  INV_X1 U30510 ( .A(n63209), .ZN(n26040) );
  INV_X1 U30511 ( .A(n26040), .ZN(p_wishbone_bd_ram_n25052) );
  INV_X1 U30512 ( .A(n63208), .ZN(n26042) );
  INV_X1 U30513 ( .A(n26042), .ZN(p_wishbone_bd_ram_n25051) );
  INV_X1 U30514 ( .A(n63207), .ZN(n26044) );
  INV_X1 U30515 ( .A(n26044), .ZN(p_wishbone_bd_ram_n25050) );
  INV_X1 U30516 ( .A(n63206), .ZN(n26046) );
  INV_X1 U30517 ( .A(n26046), .ZN(p_wishbone_bd_ram_n25049) );
  INV_X1 U30518 ( .A(n63205), .ZN(n26048) );
  INV_X1 U30519 ( .A(n26048), .ZN(p_wishbone_bd_ram_n25048) );
  INV_X1 U30520 ( .A(n63204), .ZN(n26050) );
  INV_X1 U30521 ( .A(n26050), .ZN(p_wishbone_bd_ram_n25047) );
  INV_X1 U30522 ( .A(n63203), .ZN(n26052) );
  INV_X1 U30523 ( .A(n26052), .ZN(p_wishbone_bd_ram_n25046) );
  INV_X1 U30524 ( .A(n63202), .ZN(n26054) );
  INV_X1 U30525 ( .A(n26054), .ZN(p_wishbone_bd_ram_n25045) );
  INV_X1 U30526 ( .A(n63201), .ZN(n26056) );
  INV_X1 U30527 ( .A(n26056), .ZN(p_wishbone_bd_ram_n25044) );
  INV_X1 U30528 ( .A(n63200), .ZN(n26058) );
  INV_X1 U30529 ( .A(n26058), .ZN(p_wishbone_bd_ram_n25043) );
  INV_X1 U30530 ( .A(n63199), .ZN(n26060) );
  INV_X1 U30531 ( .A(n26060), .ZN(p_wishbone_bd_ram_n25042) );
  INV_X1 U30532 ( .A(n63198), .ZN(n26062) );
  INV_X1 U30533 ( .A(n26062), .ZN(p_wishbone_bd_ram_n25041) );
  INV_X1 U30534 ( .A(n63197), .ZN(n26064) );
  INV_X1 U30535 ( .A(n26064), .ZN(p_wishbone_bd_ram_n25040) );
  INV_X1 U30536 ( .A(n63196), .ZN(n26066) );
  INV_X1 U30537 ( .A(n26066), .ZN(p_wishbone_bd_ram_n25039) );
  INV_X1 U30538 ( .A(n63195), .ZN(n26068) );
  INV_X1 U30539 ( .A(n26068), .ZN(p_wishbone_bd_ram_n25038) );
  INV_X1 U30540 ( .A(n63194), .ZN(n26070) );
  INV_X1 U30541 ( .A(n26070), .ZN(p_wishbone_bd_ram_n25037) );
  INV_X1 U30542 ( .A(n63193), .ZN(n26072) );
  INV_X1 U30543 ( .A(n26072), .ZN(p_wishbone_bd_ram_n25036) );
  INV_X1 U30544 ( .A(n63192), .ZN(n26074) );
  INV_X1 U30545 ( .A(n26074), .ZN(p_wishbone_bd_ram_n25035) );
  INV_X1 U30546 ( .A(n63191), .ZN(n26076) );
  INV_X1 U30547 ( .A(n26076), .ZN(p_wishbone_bd_ram_n25034) );
  INV_X1 U30548 ( .A(n63190), .ZN(n26078) );
  INV_X1 U30549 ( .A(n26078), .ZN(p_wishbone_bd_ram_n25033) );
  INV_X1 U30550 ( .A(n63189), .ZN(n26080) );
  INV_X1 U30551 ( .A(n26080), .ZN(p_wishbone_bd_ram_n25032) );
  INV_X1 U30552 ( .A(n63188), .ZN(n26082) );
  INV_X1 U30553 ( .A(n26082), .ZN(p_wishbone_bd_ram_n25031) );
  INV_X1 U30554 ( .A(n63187), .ZN(n26084) );
  INV_X1 U30555 ( .A(n26084), .ZN(p_wishbone_bd_ram_n25030) );
  INV_X1 U30556 ( .A(n63186), .ZN(n26086) );
  INV_X1 U30557 ( .A(n26086), .ZN(p_wishbone_bd_ram_n25029) );
  INV_X1 U30558 ( .A(n63185), .ZN(n26088) );
  INV_X1 U30559 ( .A(n26088), .ZN(p_wishbone_bd_ram_n25028) );
  INV_X1 U30560 ( .A(n63184), .ZN(n26090) );
  INV_X1 U30561 ( .A(n26090), .ZN(p_wishbone_bd_ram_n25027) );
  INV_X1 U30562 ( .A(n63183), .ZN(n26092) );
  INV_X1 U30563 ( .A(n26092), .ZN(p_wishbone_bd_ram_n25026) );
  INV_X1 U30564 ( .A(n63182), .ZN(n26094) );
  INV_X1 U30565 ( .A(n26094), .ZN(p_wishbone_bd_ram_n25025) );
  INV_X1 U30566 ( .A(n63181), .ZN(n26096) );
  INV_X1 U30567 ( .A(n26096), .ZN(p_wishbone_bd_ram_n25024) );
  INV_X1 U30568 ( .A(n63180), .ZN(n26098) );
  INV_X1 U30569 ( .A(n26098), .ZN(p_wishbone_bd_ram_n25023) );
  INV_X1 U30570 ( .A(n63179), .ZN(n26100) );
  INV_X1 U30571 ( .A(n26100), .ZN(p_wishbone_bd_ram_n25022) );
  INV_X1 U30572 ( .A(n63178), .ZN(n26102) );
  INV_X1 U30573 ( .A(n26102), .ZN(p_wishbone_bd_ram_n25021) );
  INV_X1 U30574 ( .A(n63177), .ZN(n26104) );
  INV_X1 U30575 ( .A(n26104), .ZN(p_wishbone_bd_ram_n25020) );
  INV_X1 U30576 ( .A(n63176), .ZN(n26106) );
  INV_X1 U30577 ( .A(n26106), .ZN(p_wishbone_bd_ram_n25019) );
  INV_X1 U30578 ( .A(n63175), .ZN(n26108) );
  INV_X1 U30579 ( .A(n26108), .ZN(p_wishbone_bd_ram_n25018) );
  INV_X1 U30580 ( .A(n63174), .ZN(n26110) );
  INV_X1 U30581 ( .A(n26110), .ZN(p_wishbone_bd_ram_n25017) );
  INV_X1 U30582 ( .A(n63173), .ZN(n26112) );
  INV_X1 U30583 ( .A(n26112), .ZN(p_wishbone_bd_ram_n25016) );
  INV_X1 U30584 ( .A(n63172), .ZN(n26114) );
  INV_X1 U30585 ( .A(n26114), .ZN(p_wishbone_bd_ram_n25015) );
  INV_X1 U30586 ( .A(n63171), .ZN(n26116) );
  INV_X1 U30587 ( .A(n26116), .ZN(p_wishbone_bd_ram_n25014) );
  INV_X1 U30588 ( .A(n63170), .ZN(n26118) );
  INV_X1 U30589 ( .A(n26118), .ZN(p_wishbone_bd_ram_n25013) );
  INV_X1 U30590 ( .A(n63169), .ZN(n26120) );
  INV_X1 U30591 ( .A(n26120), .ZN(p_wishbone_bd_ram_n25012) );
  INV_X1 U30592 ( .A(n63168), .ZN(n26122) );
  INV_X1 U30593 ( .A(n26122), .ZN(p_wishbone_bd_ram_n25011) );
  INV_X1 U30594 ( .A(n63167), .ZN(n26124) );
  INV_X1 U30595 ( .A(n26124), .ZN(p_wishbone_bd_ram_n25010) );
  INV_X1 U30596 ( .A(n63166), .ZN(n26126) );
  INV_X1 U30597 ( .A(n26126), .ZN(p_wishbone_bd_ram_n25009) );
  INV_X1 U30598 ( .A(n63165), .ZN(n26128) );
  INV_X1 U30599 ( .A(n26128), .ZN(p_wishbone_bd_ram_n25008) );
  INV_X1 U30600 ( .A(n63164), .ZN(n26130) );
  INV_X1 U30601 ( .A(n26130), .ZN(p_wishbone_bd_ram_n25007) );
  INV_X1 U30602 ( .A(n63163), .ZN(n26132) );
  INV_X1 U30603 ( .A(n26132), .ZN(p_wishbone_bd_ram_n25006) );
  INV_X1 U30604 ( .A(n63162), .ZN(n26134) );
  INV_X1 U30605 ( .A(n26134), .ZN(p_wishbone_bd_ram_n25005) );
  INV_X1 U30606 ( .A(n63161), .ZN(n26136) );
  INV_X1 U30607 ( .A(n26136), .ZN(p_wishbone_bd_ram_n25004) );
  INV_X1 U30608 ( .A(n63160), .ZN(n26138) );
  INV_X1 U30609 ( .A(n26138), .ZN(p_wishbone_bd_ram_n25003) );
  INV_X1 U30610 ( .A(n63159), .ZN(n26140) );
  INV_X1 U30611 ( .A(n26140), .ZN(p_wishbone_bd_ram_n25002) );
  INV_X1 U30612 ( .A(n63158), .ZN(n26142) );
  INV_X1 U30613 ( .A(n26142), .ZN(p_wishbone_bd_ram_n25001) );
  INV_X1 U30614 ( .A(n63157), .ZN(n26144) );
  INV_X1 U30615 ( .A(n26144), .ZN(p_wishbone_bd_ram_n24999) );
  INV_X1 U30616 ( .A(n63156), .ZN(n26146) );
  INV_X1 U30617 ( .A(n26146), .ZN(p_wishbone_bd_ram_n24997) );
  INV_X1 U30618 ( .A(n63155), .ZN(n26148) );
  INV_X1 U30619 ( .A(n26148), .ZN(p_wishbone_bd_ram_n24996) );
  INV_X1 U30620 ( .A(n63154), .ZN(n26150) );
  INV_X1 U30621 ( .A(n26150), .ZN(p_wishbone_bd_ram_n24994) );
  INV_X1 U30622 ( .A(n63153), .ZN(n26152) );
  INV_X1 U30623 ( .A(n26152), .ZN(p_wishbone_bd_ram_n24991) );
  INV_X1 U30624 ( .A(n63152), .ZN(n26154) );
  INV_X1 U30625 ( .A(n26154), .ZN(p_wishbone_bd_ram_n24989) );
  INV_X1 U30626 ( .A(n63151), .ZN(n26156) );
  INV_X1 U30627 ( .A(n26156), .ZN(p_wishbone_bd_ram_n24988) );
  INV_X1 U30628 ( .A(n63150), .ZN(n26158) );
  INV_X1 U30629 ( .A(n26158), .ZN(p_wishbone_bd_ram_n24986) );
  INV_X1 U30630 ( .A(n63149), .ZN(n26160) );
  INV_X1 U30631 ( .A(n26160), .ZN(p_wishbone_bd_ram_n24984) );
  INV_X1 U30632 ( .A(n63148), .ZN(n26162) );
  INV_X1 U30633 ( .A(n26162), .ZN(p_wishbone_bd_ram_n24983) );
  INV_X1 U30634 ( .A(n63147), .ZN(n26164) );
  INV_X1 U30635 ( .A(n26164), .ZN(p_wishbone_bd_ram_n24982) );
  INV_X1 U30636 ( .A(n63146), .ZN(n26166) );
  INV_X1 U30637 ( .A(n26166), .ZN(p_wishbone_bd_ram_n24981) );
  INV_X1 U30638 ( .A(n63145), .ZN(n26168) );
  INV_X1 U30639 ( .A(n26168), .ZN(p_wishbone_bd_ram_n24980) );
  INV_X1 U30640 ( .A(n63144), .ZN(n26170) );
  INV_X1 U30641 ( .A(n26170), .ZN(p_wishbone_bd_ram_n24979) );
  INV_X1 U30642 ( .A(n63143), .ZN(n26172) );
  INV_X1 U30643 ( .A(n26172), .ZN(p_wishbone_bd_ram_n24978) );
  INV_X1 U30644 ( .A(n63142), .ZN(n26174) );
  INV_X1 U30645 ( .A(n26174), .ZN(p_wishbone_bd_ram_n24977) );
  INV_X1 U30646 ( .A(n63141), .ZN(n26176) );
  INV_X1 U30647 ( .A(n26176), .ZN(p_wishbone_bd_ram_n24976) );
  INV_X1 U30648 ( .A(n63140), .ZN(n26178) );
  INV_X1 U30649 ( .A(n26178), .ZN(p_wishbone_bd_ram_n24975) );
  INV_X1 U30650 ( .A(n63139), .ZN(n26180) );
  INV_X1 U30651 ( .A(n26180), .ZN(p_wishbone_bd_ram_n24974) );
  INV_X1 U30652 ( .A(n63138), .ZN(n26182) );
  INV_X1 U30653 ( .A(n26182), .ZN(p_wishbone_bd_ram_n24973) );
  INV_X1 U30654 ( .A(n63137), .ZN(n26184) );
  INV_X1 U30655 ( .A(n26184), .ZN(p_wishbone_bd_ram_n24972) );
  INV_X1 U30656 ( .A(n63136), .ZN(n26186) );
  INV_X1 U30657 ( .A(n26186), .ZN(p_wishbone_bd_ram_n24971) );
  INV_X1 U30658 ( .A(n63135), .ZN(n26188) );
  INV_X1 U30659 ( .A(n26188), .ZN(p_wishbone_bd_ram_n24970) );
  INV_X1 U30660 ( .A(n63134), .ZN(n26190) );
  INV_X1 U30661 ( .A(n26190), .ZN(p_wishbone_bd_ram_n24969) );
  INV_X1 U30662 ( .A(n63133), .ZN(n26192) );
  INV_X1 U30663 ( .A(n26192), .ZN(p_wishbone_bd_ram_n24967) );
  INV_X1 U30664 ( .A(n63132), .ZN(n26194) );
  INV_X1 U30665 ( .A(n26194), .ZN(p_wishbone_bd_ram_n24965) );
  INV_X1 U30666 ( .A(n63131), .ZN(n26196) );
  INV_X1 U30667 ( .A(n26196), .ZN(p_wishbone_bd_ram_n24964) );
  INV_X1 U30668 ( .A(n63130), .ZN(n26198) );
  INV_X1 U30669 ( .A(n26198), .ZN(p_wishbone_bd_ram_n24962) );
  INV_X1 U30670 ( .A(n63129), .ZN(n26200) );
  INV_X1 U30671 ( .A(n26200), .ZN(p_wishbone_bd_ram_n24960) );
  INV_X1 U30672 ( .A(n63128), .ZN(n26202) );
  INV_X1 U30673 ( .A(n26202), .ZN(p_wishbone_bd_ram_n24959) );
  INV_X1 U30674 ( .A(n63127), .ZN(n26204) );
  INV_X1 U30675 ( .A(n26204), .ZN(p_wishbone_bd_ram_n24958) );
  INV_X1 U30676 ( .A(n63126), .ZN(n26206) );
  INV_X1 U30677 ( .A(n26206), .ZN(p_wishbone_bd_ram_n24957) );
  INV_X1 U30678 ( .A(n63125), .ZN(n26208) );
  INV_X1 U30679 ( .A(n26208), .ZN(p_wishbone_bd_ram_n24956) );
  INV_X1 U30680 ( .A(n63124), .ZN(n26210) );
  INV_X1 U30681 ( .A(n26210), .ZN(p_wishbone_bd_ram_n24955) );
  INV_X1 U30682 ( .A(n63123), .ZN(n26212) );
  INV_X1 U30683 ( .A(n26212), .ZN(p_wishbone_bd_ram_n24954) );
  INV_X1 U30684 ( .A(n63122), .ZN(n26214) );
  INV_X1 U30685 ( .A(n26214), .ZN(p_wishbone_bd_ram_n24953) );
  INV_X1 U30686 ( .A(n63121), .ZN(n26216) );
  INV_X1 U30687 ( .A(n26216), .ZN(p_wishbone_bd_ram_n24952) );
  INV_X1 U30688 ( .A(n63120), .ZN(n26218) );
  INV_X1 U30689 ( .A(n26218), .ZN(p_wishbone_bd_ram_n24951) );
  INV_X1 U30690 ( .A(n63119), .ZN(n26220) );
  INV_X1 U30691 ( .A(n26220), .ZN(p_wishbone_bd_ram_n24950) );
  INV_X1 U30692 ( .A(n63118), .ZN(n26222) );
  INV_X1 U30693 ( .A(n26222), .ZN(p_wishbone_bd_ram_n24949) );
  INV_X1 U30694 ( .A(n63117), .ZN(n26224) );
  INV_X1 U30695 ( .A(n26224), .ZN(p_wishbone_bd_ram_n24948) );
  INV_X1 U30696 ( .A(n63116), .ZN(n26226) );
  INV_X1 U30697 ( .A(n26226), .ZN(p_wishbone_bd_ram_n24947) );
  INV_X1 U30698 ( .A(n63115), .ZN(n26228) );
  INV_X1 U30699 ( .A(n26228), .ZN(p_wishbone_bd_ram_n24946) );
  INV_X1 U30700 ( .A(n63114), .ZN(n26230) );
  INV_X1 U30701 ( .A(n26230), .ZN(p_wishbone_bd_ram_n24945) );
  INV_X1 U30702 ( .A(n63113), .ZN(n26232) );
  INV_X1 U30703 ( .A(n26232), .ZN(p_wishbone_bd_ram_n24944) );
  INV_X1 U30704 ( .A(n63112), .ZN(n26234) );
  INV_X1 U30705 ( .A(n26234), .ZN(p_wishbone_bd_ram_n24943) );
  INV_X1 U30706 ( .A(n63111), .ZN(n26236) );
  INV_X1 U30707 ( .A(n26236), .ZN(p_wishbone_bd_ram_n24942) );
  INV_X1 U30708 ( .A(n63110), .ZN(n26238) );
  INV_X1 U30709 ( .A(n26238), .ZN(p_wishbone_bd_ram_n24941) );
  INV_X1 U30710 ( .A(n63109), .ZN(n26240) );
  INV_X1 U30711 ( .A(n26240), .ZN(p_wishbone_bd_ram_n24940) );
  INV_X1 U30712 ( .A(n63108), .ZN(n26242) );
  INV_X1 U30713 ( .A(n26242), .ZN(p_wishbone_bd_ram_n24939) );
  INV_X1 U30714 ( .A(n63107), .ZN(n26244) );
  INV_X1 U30715 ( .A(n26244), .ZN(p_wishbone_bd_ram_n24938) );
  INV_X1 U30716 ( .A(n63106), .ZN(n26246) );
  INV_X1 U30717 ( .A(n26246), .ZN(p_wishbone_bd_ram_n24937) );
  INV_X1 U30718 ( .A(n63105), .ZN(n26248) );
  INV_X1 U30719 ( .A(n26248), .ZN(p_wishbone_bd_ram_n24936) );
  INV_X1 U30720 ( .A(n63104), .ZN(n26250) );
  INV_X1 U30721 ( .A(n26250), .ZN(p_wishbone_bd_ram_n24935) );
  INV_X1 U30722 ( .A(n63103), .ZN(n26252) );
  INV_X1 U30723 ( .A(n26252), .ZN(p_wishbone_bd_ram_n24934) );
  INV_X1 U30724 ( .A(n63102), .ZN(n26254) );
  INV_X1 U30725 ( .A(n26254), .ZN(p_wishbone_bd_ram_n24933) );
  INV_X1 U30726 ( .A(n63101), .ZN(n26256) );
  INV_X1 U30727 ( .A(n26256), .ZN(p_wishbone_bd_ram_n24932) );
  INV_X1 U30728 ( .A(n63100), .ZN(n26258) );
  INV_X1 U30729 ( .A(n26258), .ZN(p_wishbone_bd_ram_n24931) );
  INV_X1 U30730 ( .A(n63099), .ZN(n26260) );
  INV_X1 U30731 ( .A(n26260), .ZN(p_wishbone_bd_ram_n24930) );
  INV_X1 U30732 ( .A(n63098), .ZN(n26262) );
  INV_X1 U30733 ( .A(n26262), .ZN(p_wishbone_bd_ram_n24929) );
  INV_X1 U30734 ( .A(n63097), .ZN(n26264) );
  INV_X1 U30735 ( .A(n26264), .ZN(p_wishbone_bd_ram_n24928) );
  INV_X1 U30736 ( .A(n63096), .ZN(n26266) );
  INV_X1 U30737 ( .A(n26266), .ZN(p_wishbone_bd_ram_n24927) );
  INV_X1 U30738 ( .A(n63095), .ZN(n26268) );
  INV_X1 U30739 ( .A(n26268), .ZN(p_wishbone_bd_ram_n24926) );
  INV_X1 U30740 ( .A(n63094), .ZN(n26270) );
  INV_X1 U30741 ( .A(n26270), .ZN(p_wishbone_bd_ram_n24925) );
  INV_X1 U30742 ( .A(n63093), .ZN(n26272) );
  INV_X1 U30743 ( .A(n26272), .ZN(p_wishbone_bd_ram_n24924) );
  INV_X1 U30744 ( .A(n63092), .ZN(n26274) );
  INV_X1 U30745 ( .A(n26274), .ZN(p_wishbone_bd_ram_n24923) );
  INV_X1 U30746 ( .A(n63091), .ZN(n26276) );
  INV_X1 U30747 ( .A(n26276), .ZN(p_wishbone_bd_ram_n24922) );
  INV_X1 U30748 ( .A(n63090), .ZN(n26278) );
  INV_X1 U30749 ( .A(n26278), .ZN(p_wishbone_bd_ram_n24921) );
  INV_X1 U30750 ( .A(n63089), .ZN(n26280) );
  INV_X1 U30751 ( .A(n26280), .ZN(p_wishbone_bd_ram_n24919) );
  INV_X1 U30752 ( .A(n63088), .ZN(n26282) );
  INV_X1 U30753 ( .A(n26282), .ZN(p_wishbone_bd_ram_n24917) );
  INV_X1 U30754 ( .A(n63087), .ZN(n26284) );
  INV_X1 U30755 ( .A(n26284), .ZN(p_wishbone_bd_ram_n24916) );
  INV_X1 U30756 ( .A(n63086), .ZN(n26286) );
  INV_X1 U30757 ( .A(n26286), .ZN(p_wishbone_bd_ram_n24914) );
  INV_X1 U30758 ( .A(n63085), .ZN(n26288) );
  INV_X1 U30759 ( .A(n26288), .ZN(p_wishbone_bd_ram_n24912) );
  INV_X1 U30760 ( .A(n63084), .ZN(n26290) );
  INV_X1 U30761 ( .A(n26290), .ZN(p_wishbone_bd_ram_n24911) );
  INV_X1 U30762 ( .A(n63083), .ZN(n26292) );
  INV_X1 U30763 ( .A(n26292), .ZN(p_wishbone_bd_ram_n24910) );
  INV_X1 U30764 ( .A(n63082), .ZN(n26294) );
  INV_X1 U30765 ( .A(n26294), .ZN(p_wishbone_bd_ram_n24909) );
  INV_X1 U30766 ( .A(n63081), .ZN(n26296) );
  INV_X1 U30767 ( .A(n26296), .ZN(p_wishbone_bd_ram_n24908) );
  INV_X1 U30768 ( .A(n63080), .ZN(n26298) );
  INV_X1 U30769 ( .A(n26298), .ZN(p_wishbone_bd_ram_n24907) );
  INV_X1 U30770 ( .A(n63079), .ZN(n26300) );
  INV_X1 U30771 ( .A(n26300), .ZN(p_wishbone_bd_ram_n24906) );
  INV_X1 U30772 ( .A(n63078), .ZN(n26302) );
  INV_X1 U30773 ( .A(n26302), .ZN(p_wishbone_bd_ram_n24905) );
  INV_X1 U30774 ( .A(n63077), .ZN(n26304) );
  INV_X1 U30775 ( .A(n26304), .ZN(p_wishbone_bd_ram_n24904) );
  INV_X1 U30776 ( .A(n63076), .ZN(n26306) );
  INV_X1 U30777 ( .A(n26306), .ZN(p_wishbone_bd_ram_n24903) );
  INV_X1 U30778 ( .A(n63075), .ZN(n26308) );
  INV_X1 U30779 ( .A(n26308), .ZN(p_wishbone_bd_ram_n24902) );
  INV_X1 U30780 ( .A(n63074), .ZN(n26310) );
  INV_X1 U30781 ( .A(n26310), .ZN(p_wishbone_bd_ram_n24901) );
  INV_X1 U30782 ( .A(n63073), .ZN(n26312) );
  INV_X1 U30783 ( .A(n26312), .ZN(p_wishbone_bd_ram_n24900) );
  INV_X1 U30784 ( .A(n63072), .ZN(n26314) );
  INV_X1 U30785 ( .A(n26314), .ZN(p_wishbone_bd_ram_n24899) );
  INV_X1 U30786 ( .A(n63071), .ZN(n26316) );
  INV_X1 U30787 ( .A(n26316), .ZN(p_wishbone_bd_ram_n24898) );
  INV_X1 U30788 ( .A(n63070), .ZN(n26318) );
  INV_X1 U30789 ( .A(n26318), .ZN(p_wishbone_bd_ram_n24897) );
  INV_X1 U30790 ( .A(n63069), .ZN(n26320) );
  INV_X1 U30791 ( .A(n26320), .ZN(p_wishbone_bd_ram_n24895) );
  INV_X1 U30792 ( .A(n63068), .ZN(n26322) );
  INV_X1 U30793 ( .A(n26322), .ZN(p_wishbone_bd_ram_n24893) );
  INV_X1 U30794 ( .A(n63067), .ZN(n26324) );
  INV_X1 U30795 ( .A(n26324), .ZN(p_wishbone_bd_ram_n24892) );
  INV_X1 U30796 ( .A(n63066), .ZN(n26326) );
  INV_X1 U30797 ( .A(n26326), .ZN(p_wishbone_bd_ram_n24890) );
  INV_X1 U30798 ( .A(n63065), .ZN(n26328) );
  INV_X1 U30799 ( .A(n26328), .ZN(p_wishbone_bd_ram_n24888) );
  INV_X1 U30800 ( .A(n63064), .ZN(n26330) );
  INV_X1 U30801 ( .A(n26330), .ZN(p_wishbone_bd_ram_n24887) );
  INV_X1 U30802 ( .A(n63063), .ZN(n26332) );
  INV_X1 U30803 ( .A(n26332), .ZN(p_wishbone_bd_ram_n24886) );
  INV_X1 U30804 ( .A(n63062), .ZN(n26334) );
  INV_X1 U30805 ( .A(n26334), .ZN(p_wishbone_bd_ram_n24885) );
  INV_X1 U30806 ( .A(n63061), .ZN(n26336) );
  INV_X1 U30807 ( .A(n26336), .ZN(p_wishbone_bd_ram_n24884) );
  INV_X1 U30808 ( .A(n63060), .ZN(n26338) );
  INV_X1 U30809 ( .A(n26338), .ZN(p_wishbone_bd_ram_n24883) );
  INV_X1 U30810 ( .A(n63059), .ZN(n26340) );
  INV_X1 U30811 ( .A(n26340), .ZN(p_wishbone_bd_ram_n24882) );
  INV_X1 U30812 ( .A(n63058), .ZN(n26342) );
  INV_X1 U30813 ( .A(n26342), .ZN(p_wishbone_bd_ram_n24881) );
  INV_X1 U30814 ( .A(n63057), .ZN(n26344) );
  INV_X1 U30815 ( .A(n26344), .ZN(p_wishbone_bd_ram_n24880) );
  INV_X1 U30816 ( .A(n63056), .ZN(n26346) );
  INV_X1 U30817 ( .A(n26346), .ZN(p_wishbone_bd_ram_n24879) );
  INV_X1 U30818 ( .A(n63055), .ZN(n26348) );
  INV_X1 U30819 ( .A(n26348), .ZN(p_wishbone_bd_ram_n24878) );
  INV_X1 U30820 ( .A(n63054), .ZN(n26350) );
  INV_X1 U30821 ( .A(n26350), .ZN(p_wishbone_bd_ram_n24877) );
  INV_X1 U30822 ( .A(n63053), .ZN(n26352) );
  INV_X1 U30823 ( .A(n26352), .ZN(p_wishbone_bd_ram_n24876) );
  INV_X1 U30824 ( .A(n63052), .ZN(n26354) );
  INV_X1 U30825 ( .A(n26354), .ZN(p_wishbone_bd_ram_n24875) );
  INV_X1 U30826 ( .A(n63051), .ZN(n26356) );
  INV_X1 U30827 ( .A(n26356), .ZN(p_wishbone_bd_ram_n24874) );
  INV_X1 U30828 ( .A(n63050), .ZN(n26358) );
  INV_X1 U30829 ( .A(n26358), .ZN(p_wishbone_bd_ram_n24873) );
  INV_X1 U30830 ( .A(n63049), .ZN(n26360) );
  INV_X1 U30831 ( .A(n26360), .ZN(p_wishbone_bd_ram_n24872) );
  INV_X1 U30832 ( .A(n63048), .ZN(n26362) );
  INV_X1 U30833 ( .A(n26362), .ZN(p_wishbone_bd_ram_n24871) );
  INV_X1 U30834 ( .A(n63047), .ZN(n26364) );
  INV_X1 U30835 ( .A(n26364), .ZN(p_wishbone_bd_ram_n24870) );
  INV_X1 U30836 ( .A(n63046), .ZN(n26366) );
  INV_X1 U30837 ( .A(n26366), .ZN(p_wishbone_bd_ram_n24869) );
  INV_X1 U30838 ( .A(n63045), .ZN(n26368) );
  INV_X1 U30839 ( .A(n26368), .ZN(p_wishbone_bd_ram_n24868) );
  INV_X1 U30840 ( .A(n63044), .ZN(n26370) );
  INV_X1 U30841 ( .A(n26370), .ZN(p_wishbone_bd_ram_n24867) );
  INV_X1 U30842 ( .A(n63043), .ZN(n26372) );
  INV_X1 U30843 ( .A(n26372), .ZN(p_wishbone_bd_ram_n24866) );
  INV_X1 U30844 ( .A(n63042), .ZN(n26374) );
  INV_X1 U30845 ( .A(n26374), .ZN(p_wishbone_bd_ram_n24865) );
  INV_X1 U30846 ( .A(n63041), .ZN(n26376) );
  INV_X1 U30847 ( .A(n26376), .ZN(p_wishbone_bd_ram_n24864) );
  INV_X1 U30848 ( .A(n63040), .ZN(n26378) );
  INV_X1 U30849 ( .A(n26378), .ZN(p_wishbone_bd_ram_n24863) );
  INV_X1 U30850 ( .A(n63039), .ZN(n26380) );
  INV_X1 U30851 ( .A(n26380), .ZN(p_wishbone_bd_ram_n24862) );
  INV_X1 U30852 ( .A(n63038), .ZN(n26382) );
  INV_X1 U30853 ( .A(n26382), .ZN(p_wishbone_bd_ram_n24861) );
  INV_X1 U30854 ( .A(n63037), .ZN(n26384) );
  INV_X1 U30855 ( .A(n26384), .ZN(p_wishbone_bd_ram_n24860) );
  INV_X1 U30856 ( .A(n63036), .ZN(n26386) );
  INV_X1 U30857 ( .A(n26386), .ZN(p_wishbone_bd_ram_n24859) );
  INV_X1 U30858 ( .A(n63035), .ZN(n26388) );
  INV_X1 U30859 ( .A(n26388), .ZN(p_wishbone_bd_ram_n24858) );
  INV_X1 U30860 ( .A(n63034), .ZN(n26390) );
  INV_X1 U30861 ( .A(n26390), .ZN(p_wishbone_bd_ram_n24857) );
  INV_X1 U30862 ( .A(n63033), .ZN(n26392) );
  INV_X1 U30863 ( .A(n26392), .ZN(p_wishbone_bd_ram_n24856) );
  INV_X1 U30864 ( .A(n63032), .ZN(n26394) );
  INV_X1 U30865 ( .A(n26394), .ZN(p_wishbone_bd_ram_n24855) );
  INV_X1 U30866 ( .A(n63031), .ZN(n26396) );
  INV_X1 U30867 ( .A(n26396), .ZN(p_wishbone_bd_ram_n24854) );
  INV_X1 U30868 ( .A(n63030), .ZN(n26398) );
  INV_X1 U30869 ( .A(n26398), .ZN(p_wishbone_bd_ram_n24853) );
  INV_X1 U30870 ( .A(n63029), .ZN(n26400) );
  INV_X1 U30871 ( .A(n26400), .ZN(p_wishbone_bd_ram_n24852) );
  INV_X1 U30872 ( .A(n63028), .ZN(n26402) );
  INV_X1 U30873 ( .A(n26402), .ZN(p_wishbone_bd_ram_n24851) );
  INV_X1 U30874 ( .A(n63027), .ZN(n26404) );
  INV_X1 U30875 ( .A(n26404), .ZN(p_wishbone_bd_ram_n24850) );
  INV_X1 U30876 ( .A(n63026), .ZN(n26406) );
  INV_X1 U30877 ( .A(n26406), .ZN(p_wishbone_bd_ram_n24849) );
  INV_X1 U30878 ( .A(n63025), .ZN(n26408) );
  INV_X1 U30879 ( .A(n26408), .ZN(p_wishbone_bd_ram_n24848) );
  INV_X1 U30880 ( .A(n63024), .ZN(n26410) );
  INV_X1 U30881 ( .A(n26410), .ZN(p_wishbone_bd_ram_n24847) );
  INV_X1 U30882 ( .A(n63023), .ZN(n26412) );
  INV_X1 U30883 ( .A(n26412), .ZN(p_wishbone_bd_ram_n24846) );
  INV_X1 U30884 ( .A(n63022), .ZN(n26414) );
  INV_X1 U30885 ( .A(n26414), .ZN(p_wishbone_bd_ram_n24845) );
  INV_X1 U30886 ( .A(n63021), .ZN(n26416) );
  INV_X1 U30887 ( .A(n26416), .ZN(p_wishbone_bd_ram_n24844) );
  INV_X1 U30888 ( .A(n63020), .ZN(n26418) );
  INV_X1 U30889 ( .A(n26418), .ZN(p_wishbone_bd_ram_n24843) );
  INV_X1 U30890 ( .A(n63019), .ZN(n26420) );
  INV_X1 U30891 ( .A(n26420), .ZN(p_wishbone_bd_ram_n24842) );
  INV_X1 U30892 ( .A(n63018), .ZN(n26422) );
  INV_X1 U30893 ( .A(n26422), .ZN(p_wishbone_bd_ram_n24841) );
  INV_X1 U30894 ( .A(n63017), .ZN(n26424) );
  INV_X1 U30895 ( .A(n26424), .ZN(p_wishbone_bd_ram_n24840) );
  INV_X1 U30896 ( .A(n63016), .ZN(n26426) );
  INV_X1 U30897 ( .A(n26426), .ZN(p_wishbone_bd_ram_n24839) );
  INV_X1 U30898 ( .A(n63015), .ZN(n26428) );
  INV_X1 U30899 ( .A(n26428), .ZN(p_wishbone_bd_ram_n24838) );
  INV_X1 U30900 ( .A(n63014), .ZN(n26430) );
  INV_X1 U30901 ( .A(n26430), .ZN(p_wishbone_bd_ram_n24837) );
  INV_X1 U30902 ( .A(n63013), .ZN(n26432) );
  INV_X1 U30903 ( .A(n26432), .ZN(p_wishbone_bd_ram_n24836) );
  INV_X1 U30904 ( .A(n63012), .ZN(n26434) );
  INV_X1 U30905 ( .A(n26434), .ZN(p_wishbone_bd_ram_n24835) );
  INV_X1 U30906 ( .A(n63011), .ZN(n26436) );
  INV_X1 U30907 ( .A(n26436), .ZN(p_wishbone_bd_ram_n24834) );
  INV_X1 U30908 ( .A(n63010), .ZN(n26438) );
  INV_X1 U30909 ( .A(n26438), .ZN(p_wishbone_bd_ram_n24833) );
  INV_X1 U30910 ( .A(n63009), .ZN(n26440) );
  INV_X1 U30911 ( .A(n26440), .ZN(p_wishbone_bd_ram_n24831) );
  INV_X1 U30912 ( .A(n63008), .ZN(n26442) );
  INV_X1 U30913 ( .A(n26442), .ZN(p_wishbone_bd_ram_n24829) );
  INV_X1 U30914 ( .A(n63007), .ZN(n26444) );
  INV_X1 U30915 ( .A(n26444), .ZN(p_wishbone_bd_ram_n24828) );
  INV_X1 U30916 ( .A(n63006), .ZN(n26446) );
  INV_X1 U30917 ( .A(n26446), .ZN(p_wishbone_bd_ram_n24826) );
  INV_X1 U30918 ( .A(n63005), .ZN(n26448) );
  INV_X1 U30919 ( .A(n26448), .ZN(p_wishbone_bd_ram_n24823) );
  INV_X1 U30920 ( .A(n63004), .ZN(n26450) );
  INV_X1 U30921 ( .A(n26450), .ZN(p_wishbone_bd_ram_n24821) );
  INV_X1 U30922 ( .A(n63003), .ZN(n26452) );
  INV_X1 U30923 ( .A(n26452), .ZN(p_wishbone_bd_ram_n24820) );
  INV_X1 U30924 ( .A(n63002), .ZN(n26454) );
  INV_X1 U30925 ( .A(n26454), .ZN(p_wishbone_bd_ram_n24818) );
  INV_X1 U30926 ( .A(n63001), .ZN(n26456) );
  INV_X1 U30927 ( .A(n26456), .ZN(p_wishbone_bd_ram_n24816) );
  INV_X1 U30928 ( .A(n63000), .ZN(n26458) );
  INV_X1 U30929 ( .A(n26458), .ZN(p_wishbone_bd_ram_n24815) );
  INV_X1 U30930 ( .A(n62999), .ZN(n26460) );
  INV_X1 U30931 ( .A(n26460), .ZN(p_wishbone_bd_ram_n24814) );
  INV_X1 U30932 ( .A(n62998), .ZN(n26462) );
  INV_X1 U30933 ( .A(n26462), .ZN(p_wishbone_bd_ram_n24813) );
  INV_X1 U30934 ( .A(n62997), .ZN(n26464) );
  INV_X1 U30935 ( .A(n26464), .ZN(p_wishbone_bd_ram_n24812) );
  INV_X1 U30936 ( .A(n62996), .ZN(n26466) );
  INV_X1 U30937 ( .A(n26466), .ZN(p_wishbone_bd_ram_n24811) );
  INV_X1 U30938 ( .A(n62995), .ZN(n26468) );
  INV_X1 U30939 ( .A(n26468), .ZN(p_wishbone_bd_ram_n24810) );
  INV_X1 U30940 ( .A(n62994), .ZN(n26470) );
  INV_X1 U30941 ( .A(n26470), .ZN(p_wishbone_bd_ram_n24809) );
  INV_X1 U30942 ( .A(n62993), .ZN(n26472) );
  INV_X1 U30943 ( .A(n26472), .ZN(p_wishbone_bd_ram_n24807) );
  INV_X1 U30944 ( .A(n62992), .ZN(n26474) );
  INV_X1 U30945 ( .A(n26474), .ZN(p_wishbone_bd_ram_n24805) );
  INV_X1 U30946 ( .A(n62991), .ZN(n26476) );
  INV_X1 U30947 ( .A(n26476), .ZN(p_wishbone_bd_ram_n24804) );
  INV_X1 U30948 ( .A(n62990), .ZN(n26478) );
  INV_X1 U30949 ( .A(n26478), .ZN(p_wishbone_bd_ram_n24802) );
  INV_X1 U30950 ( .A(n62989), .ZN(n26480) );
  INV_X1 U30951 ( .A(n26480), .ZN(p_wishbone_bd_ram_n24800) );
  INV_X1 U30952 ( .A(n62988), .ZN(n26482) );
  INV_X1 U30953 ( .A(n26482), .ZN(p_wishbone_bd_ram_n24799) );
  INV_X1 U30954 ( .A(n62987), .ZN(n26484) );
  INV_X1 U30955 ( .A(n26484), .ZN(p_wishbone_bd_ram_n24798) );
  INV_X1 U30956 ( .A(n62986), .ZN(n26486) );
  INV_X1 U30957 ( .A(n26486), .ZN(p_wishbone_bd_ram_n24797) );
  INV_X1 U30958 ( .A(n62985), .ZN(n26488) );
  INV_X1 U30959 ( .A(n26488), .ZN(p_wishbone_bd_ram_n24796) );
  INV_X1 U30960 ( .A(n62984), .ZN(n26490) );
  INV_X1 U30961 ( .A(n26490), .ZN(p_wishbone_bd_ram_n24795) );
  INV_X1 U30962 ( .A(n62983), .ZN(n26492) );
  INV_X1 U30963 ( .A(n26492), .ZN(p_wishbone_bd_ram_n24794) );
  INV_X1 U30964 ( .A(n62982), .ZN(n26494) );
  INV_X1 U30965 ( .A(n26494), .ZN(p_wishbone_bd_ram_n24793) );
  INV_X1 U30966 ( .A(n62981), .ZN(n26496) );
  INV_X1 U30967 ( .A(n26496), .ZN(p_wishbone_bd_ram_n24792) );
  INV_X1 U30968 ( .A(n62980), .ZN(n26498) );
  INV_X1 U30969 ( .A(n26498), .ZN(p_wishbone_bd_ram_n24791) );
  INV_X1 U30970 ( .A(n62979), .ZN(n26500) );
  INV_X1 U30971 ( .A(n26500), .ZN(p_wishbone_bd_ram_n24790) );
  INV_X1 U30972 ( .A(n62978), .ZN(n26502) );
  INV_X1 U30973 ( .A(n26502), .ZN(p_wishbone_bd_ram_n24789) );
  INV_X1 U30974 ( .A(n62977), .ZN(n26504) );
  INV_X1 U30975 ( .A(n26504), .ZN(p_wishbone_bd_ram_n24788) );
  INV_X1 U30976 ( .A(n62976), .ZN(n26506) );
  INV_X1 U30977 ( .A(n26506), .ZN(p_wishbone_bd_ram_n24787) );
  INV_X1 U30978 ( .A(n62975), .ZN(n26508) );
  INV_X1 U30979 ( .A(n26508), .ZN(p_wishbone_bd_ram_n24786) );
  INV_X1 U30980 ( .A(n62974), .ZN(n26510) );
  INV_X1 U30981 ( .A(n26510), .ZN(p_wishbone_bd_ram_n24785) );
  INV_X1 U30982 ( .A(n62973), .ZN(n26512) );
  INV_X1 U30983 ( .A(n26512), .ZN(p_wishbone_bd_ram_n24784) );
  INV_X1 U30984 ( .A(n62972), .ZN(n26514) );
  INV_X1 U30985 ( .A(n26514), .ZN(p_wishbone_bd_ram_n24783) );
  INV_X1 U30986 ( .A(n62971), .ZN(n26516) );
  INV_X1 U30987 ( .A(n26516), .ZN(p_wishbone_bd_ram_n24782) );
  INV_X1 U30988 ( .A(n62970), .ZN(n26518) );
  INV_X1 U30989 ( .A(n26518), .ZN(p_wishbone_bd_ram_n24781) );
  INV_X1 U30990 ( .A(n62969), .ZN(n26520) );
  INV_X1 U30991 ( .A(n26520), .ZN(p_wishbone_bd_ram_n24780) );
  INV_X1 U30992 ( .A(n62968), .ZN(n26522) );
  INV_X1 U30993 ( .A(n26522), .ZN(p_wishbone_bd_ram_n24779) );
  INV_X1 U30994 ( .A(n62967), .ZN(n26524) );
  INV_X1 U30995 ( .A(n26524), .ZN(p_wishbone_bd_ram_n24778) );
  INV_X1 U30996 ( .A(n62966), .ZN(n26526) );
  INV_X1 U30997 ( .A(n26526), .ZN(p_wishbone_bd_ram_n24777) );
  INV_X1 U30998 ( .A(n62965), .ZN(n26528) );
  INV_X1 U30999 ( .A(n26528), .ZN(p_wishbone_bd_ram_n24776) );
  INV_X1 U31000 ( .A(n62964), .ZN(n26530) );
  INV_X1 U31001 ( .A(n26530), .ZN(p_wishbone_bd_ram_n24775) );
  INV_X1 U31002 ( .A(n62963), .ZN(n26532) );
  INV_X1 U31003 ( .A(n26532), .ZN(p_wishbone_bd_ram_n24774) );
  INV_X1 U31004 ( .A(n62962), .ZN(n26534) );
  INV_X1 U31005 ( .A(n26534), .ZN(p_wishbone_bd_ram_n24773) );
  INV_X1 U31006 ( .A(n62961), .ZN(n26536) );
  INV_X1 U31007 ( .A(n26536), .ZN(p_wishbone_bd_ram_n24772) );
  INV_X1 U31008 ( .A(n62960), .ZN(n26538) );
  INV_X1 U31009 ( .A(n26538), .ZN(p_wishbone_bd_ram_n24771) );
  INV_X1 U31010 ( .A(n62959), .ZN(n26540) );
  INV_X1 U31011 ( .A(n26540), .ZN(p_wishbone_bd_ram_n24770) );
  INV_X1 U31012 ( .A(n62958), .ZN(n26542) );
  INV_X1 U31013 ( .A(n26542), .ZN(p_wishbone_bd_ram_n24769) );
  INV_X1 U31014 ( .A(n62957), .ZN(n26544) );
  INV_X1 U31015 ( .A(n26544), .ZN(p_wishbone_bd_ram_n24767) );
  INV_X1 U31016 ( .A(n62956), .ZN(n26546) );
  INV_X1 U31017 ( .A(n26546), .ZN(p_wishbone_bd_ram_n24765) );
  INV_X1 U31018 ( .A(n62955), .ZN(n26548) );
  INV_X1 U31019 ( .A(n26548), .ZN(p_wishbone_bd_ram_n24764) );
  INV_X1 U31020 ( .A(n62954), .ZN(n26550) );
  INV_X1 U31021 ( .A(n26550), .ZN(p_wishbone_bd_ram_n24762) );
  INV_X1 U31022 ( .A(n62953), .ZN(n26552) );
  INV_X1 U31023 ( .A(n26552), .ZN(p_wishbone_bd_ram_n24760) );
  INV_X1 U31024 ( .A(n62952), .ZN(n26554) );
  INV_X1 U31025 ( .A(n26554), .ZN(p_wishbone_bd_ram_n24759) );
  INV_X1 U31026 ( .A(n62951), .ZN(n26556) );
  INV_X1 U31027 ( .A(n26556), .ZN(p_wishbone_bd_ram_n24758) );
  INV_X1 U31028 ( .A(n62950), .ZN(n26558) );
  INV_X1 U31029 ( .A(n26558), .ZN(p_wishbone_bd_ram_n24757) );
  INV_X1 U31030 ( .A(n62949), .ZN(n26560) );
  INV_X1 U31031 ( .A(n26560), .ZN(p_wishbone_bd_ram_n24756) );
  INV_X1 U31032 ( .A(n62948), .ZN(n26562) );
  INV_X1 U31033 ( .A(n26562), .ZN(p_wishbone_bd_ram_n24755) );
  INV_X1 U31034 ( .A(n62947), .ZN(n26564) );
  INV_X1 U31035 ( .A(n26564), .ZN(p_wishbone_bd_ram_n24754) );
  INV_X1 U31036 ( .A(n62946), .ZN(n26566) );
  INV_X1 U31037 ( .A(n26566), .ZN(p_wishbone_bd_ram_n24753) );
  INV_X1 U31038 ( .A(n62945), .ZN(n26568) );
  INV_X1 U31039 ( .A(n26568), .ZN(p_wishbone_bd_ram_n24752) );
  INV_X1 U31040 ( .A(n62944), .ZN(n26570) );
  INV_X1 U31041 ( .A(n26570), .ZN(p_wishbone_bd_ram_n24751) );
  INV_X1 U31042 ( .A(n62943), .ZN(n26572) );
  INV_X1 U31043 ( .A(n26572), .ZN(p_wishbone_bd_ram_n24750) );
  INV_X1 U31044 ( .A(n62942), .ZN(n26574) );
  INV_X1 U31045 ( .A(n26574), .ZN(p_wishbone_bd_ram_n24749) );
  INV_X1 U31046 ( .A(n62941), .ZN(n26576) );
  INV_X1 U31047 ( .A(n26576), .ZN(p_wishbone_bd_ram_n24748) );
  INV_X1 U31048 ( .A(n62940), .ZN(n26578) );
  INV_X1 U31049 ( .A(n26578), .ZN(p_wishbone_bd_ram_n24747) );
  INV_X1 U31050 ( .A(n62939), .ZN(n26580) );
  INV_X1 U31051 ( .A(n26580), .ZN(p_wishbone_bd_ram_n24746) );
  INV_X1 U31052 ( .A(n62938), .ZN(n26582) );
  INV_X1 U31053 ( .A(n26582), .ZN(p_wishbone_bd_ram_n24745) );
  INV_X1 U31054 ( .A(n62937), .ZN(n26584) );
  INV_X1 U31055 ( .A(n26584), .ZN(p_wishbone_bd_ram_n24744) );
  INV_X1 U31056 ( .A(n62936), .ZN(n26586) );
  INV_X1 U31057 ( .A(n26586), .ZN(p_wishbone_bd_ram_n24743) );
  INV_X1 U31058 ( .A(n62935), .ZN(n26588) );
  INV_X1 U31059 ( .A(n26588), .ZN(p_wishbone_bd_ram_n24742) );
  INV_X1 U31060 ( .A(n62934), .ZN(n26590) );
  INV_X1 U31061 ( .A(n26590), .ZN(p_wishbone_bd_ram_n24741) );
  INV_X1 U31062 ( .A(n62933), .ZN(n26592) );
  INV_X1 U31063 ( .A(n26592), .ZN(p_wishbone_bd_ram_n24740) );
  INV_X1 U31064 ( .A(n62932), .ZN(n26594) );
  INV_X1 U31065 ( .A(n26594), .ZN(p_wishbone_bd_ram_n24739) );
  INV_X1 U31066 ( .A(n62931), .ZN(n26596) );
  INV_X1 U31067 ( .A(n26596), .ZN(p_wishbone_bd_ram_n24738) );
  INV_X1 U31068 ( .A(n62930), .ZN(n26598) );
  INV_X1 U31069 ( .A(n26598), .ZN(p_wishbone_bd_ram_n24737) );
  INV_X1 U31070 ( .A(n62929), .ZN(n26600) );
  INV_X1 U31071 ( .A(n26600), .ZN(p_wishbone_bd_ram_n24736) );
  INV_X1 U31072 ( .A(n62928), .ZN(n26602) );
  INV_X1 U31073 ( .A(n26602), .ZN(p_wishbone_bd_ram_n24735) );
  INV_X1 U31074 ( .A(n62927), .ZN(n26604) );
  INV_X1 U31075 ( .A(n26604), .ZN(p_wishbone_bd_ram_n24734) );
  INV_X1 U31076 ( .A(n62926), .ZN(n26606) );
  INV_X1 U31077 ( .A(n26606), .ZN(p_wishbone_bd_ram_n24733) );
  INV_X1 U31078 ( .A(n62925), .ZN(n26608) );
  INV_X1 U31079 ( .A(n26608), .ZN(p_wishbone_bd_ram_n24732) );
  INV_X1 U31080 ( .A(n62924), .ZN(n26610) );
  INV_X1 U31081 ( .A(n26610), .ZN(p_wishbone_bd_ram_n24731) );
  INV_X1 U31082 ( .A(n62923), .ZN(n26612) );
  INV_X1 U31083 ( .A(n26612), .ZN(p_wishbone_bd_ram_n24730) );
  INV_X1 U31084 ( .A(n62922), .ZN(n26614) );
  INV_X1 U31085 ( .A(n26614), .ZN(p_wishbone_bd_ram_n24729) );
  INV_X1 U31086 ( .A(n62921), .ZN(n26616) );
  INV_X1 U31087 ( .A(n26616), .ZN(p_wishbone_bd_ram_n24728) );
  INV_X1 U31088 ( .A(n62920), .ZN(n26618) );
  INV_X1 U31089 ( .A(n26618), .ZN(p_wishbone_bd_ram_n24727) );
  INV_X1 U31090 ( .A(n62919), .ZN(n26620) );
  INV_X1 U31091 ( .A(n26620), .ZN(p_wishbone_bd_ram_n24726) );
  INV_X1 U31092 ( .A(n62918), .ZN(n26622) );
  INV_X1 U31093 ( .A(n26622), .ZN(p_wishbone_bd_ram_n24725) );
  INV_X1 U31094 ( .A(n62917), .ZN(n26624) );
  INV_X1 U31095 ( .A(n26624), .ZN(p_wishbone_bd_ram_n24724) );
  INV_X1 U31096 ( .A(n62916), .ZN(n26626) );
  INV_X1 U31097 ( .A(n26626), .ZN(p_wishbone_bd_ram_n24723) );
  INV_X1 U31098 ( .A(n62915), .ZN(n26628) );
  INV_X1 U31099 ( .A(n26628), .ZN(p_wishbone_bd_ram_n24722) );
  INV_X1 U31100 ( .A(n62914), .ZN(n26630) );
  INV_X1 U31101 ( .A(n26630), .ZN(p_wishbone_bd_ram_n24721) );
  INV_X1 U31102 ( .A(n62913), .ZN(n26632) );
  INV_X1 U31103 ( .A(n26632), .ZN(p_wishbone_bd_ram_n24720) );
  INV_X1 U31104 ( .A(n62912), .ZN(n26634) );
  INV_X1 U31105 ( .A(n26634), .ZN(p_wishbone_bd_ram_n24719) );
  INV_X1 U31106 ( .A(n62911), .ZN(n26636) );
  INV_X1 U31107 ( .A(n26636), .ZN(p_wishbone_bd_ram_n24718) );
  INV_X1 U31108 ( .A(n62910), .ZN(n26638) );
  INV_X1 U31109 ( .A(n26638), .ZN(p_wishbone_bd_ram_n24717) );
  INV_X1 U31110 ( .A(n62909), .ZN(n26640) );
  INV_X1 U31111 ( .A(n26640), .ZN(p_wishbone_bd_ram_n24716) );
  INV_X1 U31112 ( .A(n62908), .ZN(n26642) );
  INV_X1 U31113 ( .A(n26642), .ZN(p_wishbone_bd_ram_n24715) );
  INV_X1 U31114 ( .A(n62907), .ZN(n26644) );
  INV_X1 U31115 ( .A(n26644), .ZN(p_wishbone_bd_ram_n24714) );
  INV_X1 U31116 ( .A(n62906), .ZN(n26646) );
  INV_X1 U31117 ( .A(n26646), .ZN(p_wishbone_bd_ram_n24713) );
  INV_X1 U31118 ( .A(n62905), .ZN(n26648) );
  INV_X1 U31119 ( .A(n26648), .ZN(p_wishbone_bd_ram_n24712) );
  INV_X1 U31120 ( .A(n62904), .ZN(n26650) );
  INV_X1 U31121 ( .A(n26650), .ZN(p_wishbone_bd_ram_n24711) );
  INV_X1 U31122 ( .A(n62903), .ZN(n26652) );
  INV_X1 U31123 ( .A(n26652), .ZN(p_wishbone_bd_ram_n24710) );
  INV_X1 U31124 ( .A(n62902), .ZN(n26654) );
  INV_X1 U31125 ( .A(n26654), .ZN(p_wishbone_bd_ram_n24709) );
  INV_X1 U31126 ( .A(n62901), .ZN(n26656) );
  INV_X1 U31127 ( .A(n26656), .ZN(p_wishbone_bd_ram_n24708) );
  INV_X1 U31128 ( .A(n62900), .ZN(n26658) );
  INV_X1 U31129 ( .A(n26658), .ZN(p_wishbone_bd_ram_n24707) );
  INV_X1 U31130 ( .A(n62899), .ZN(n26660) );
  INV_X1 U31131 ( .A(n26660), .ZN(p_wishbone_bd_ram_n24706) );
  INV_X1 U31132 ( .A(n62898), .ZN(n26662) );
  INV_X1 U31133 ( .A(n26662), .ZN(p_wishbone_bd_ram_n24705) );
  INV_X1 U31134 ( .A(n62897), .ZN(n26664) );
  INV_X1 U31135 ( .A(n26664), .ZN(p_wishbone_bd_ram_n24703) );
  INV_X1 U31136 ( .A(n62896), .ZN(n26666) );
  INV_X1 U31137 ( .A(n26666), .ZN(p_wishbone_bd_ram_n24701) );
  INV_X1 U31138 ( .A(n62895), .ZN(n26668) );
  INV_X1 U31139 ( .A(n26668), .ZN(p_wishbone_bd_ram_n24700) );
  INV_X1 U31140 ( .A(n62894), .ZN(n26670) );
  INV_X1 U31141 ( .A(n26670), .ZN(p_wishbone_bd_ram_n24698) );
  INV_X1 U31142 ( .A(n62893), .ZN(n26672) );
  INV_X1 U31143 ( .A(n26672), .ZN(p_wishbone_bd_ram_n24696) );
  INV_X1 U31144 ( .A(n62892), .ZN(n26674) );
  INV_X1 U31145 ( .A(n26674), .ZN(p_wishbone_bd_ram_n24695) );
  INV_X1 U31146 ( .A(n62891), .ZN(n26676) );
  INV_X1 U31147 ( .A(n26676), .ZN(p_wishbone_bd_ram_n24694) );
  INV_X1 U31148 ( .A(n62890), .ZN(n26678) );
  INV_X1 U31149 ( .A(n26678), .ZN(p_wishbone_bd_ram_n24693) );
  INV_X1 U31150 ( .A(n62889), .ZN(n26680) );
  INV_X1 U31151 ( .A(n26680), .ZN(p_wishbone_bd_ram_n24692) );
  INV_X1 U31152 ( .A(n62888), .ZN(n26682) );
  INV_X1 U31153 ( .A(n26682), .ZN(p_wishbone_bd_ram_n24691) );
  INV_X1 U31154 ( .A(n62887), .ZN(n26684) );
  INV_X1 U31155 ( .A(n26684), .ZN(p_wishbone_bd_ram_n24690) );
  INV_X1 U31156 ( .A(n62886), .ZN(n26686) );
  INV_X1 U31157 ( .A(n26686), .ZN(p_wishbone_bd_ram_n24689) );
  INV_X1 U31158 ( .A(n62885), .ZN(n26688) );
  INV_X1 U31159 ( .A(n26688), .ZN(p_wishbone_bd_ram_n24688) );
  INV_X1 U31160 ( .A(n62884), .ZN(n26690) );
  INV_X1 U31161 ( .A(n26690), .ZN(p_wishbone_bd_ram_n24687) );
  INV_X1 U31162 ( .A(n62883), .ZN(n26692) );
  INV_X1 U31163 ( .A(n26692), .ZN(p_wishbone_bd_ram_n24686) );
  INV_X1 U31164 ( .A(n62882), .ZN(n26694) );
  INV_X1 U31165 ( .A(n26694), .ZN(p_wishbone_bd_ram_n24685) );
  INV_X1 U31166 ( .A(n62881), .ZN(n26696) );
  INV_X1 U31167 ( .A(n26696), .ZN(p_wishbone_bd_ram_n24684) );
  INV_X1 U31168 ( .A(n62880), .ZN(n26698) );
  INV_X1 U31169 ( .A(n26698), .ZN(p_wishbone_bd_ram_n24683) );
  INV_X1 U31170 ( .A(n62879), .ZN(n26700) );
  INV_X1 U31171 ( .A(n26700), .ZN(p_wishbone_bd_ram_n24682) );
  INV_X1 U31172 ( .A(n62878), .ZN(n26702) );
  INV_X1 U31173 ( .A(n26702), .ZN(p_wishbone_bd_ram_n24681) );
  INV_X1 U31174 ( .A(n62877), .ZN(n26704) );
  INV_X1 U31175 ( .A(n26704), .ZN(p_wishbone_bd_ram_n24679) );
  INV_X1 U31176 ( .A(n62876), .ZN(n26706) );
  INV_X1 U31177 ( .A(n26706), .ZN(p_wishbone_bd_ram_n24677) );
  INV_X1 U31178 ( .A(n62875), .ZN(n26708) );
  INV_X1 U31179 ( .A(n26708), .ZN(p_wishbone_bd_ram_n24676) );
  INV_X1 U31180 ( .A(n62874), .ZN(n26710) );
  INV_X1 U31181 ( .A(n26710), .ZN(p_wishbone_bd_ram_n24674) );
  INV_X1 U31182 ( .A(n62873), .ZN(n26712) );
  INV_X1 U31183 ( .A(n26712), .ZN(p_wishbone_bd_ram_n24672) );
  INV_X1 U31184 ( .A(n62872), .ZN(n26714) );
  INV_X1 U31185 ( .A(n26714), .ZN(p_wishbone_bd_ram_n24671) );
  INV_X1 U31186 ( .A(n62871), .ZN(n26716) );
  INV_X1 U31187 ( .A(n26716), .ZN(p_wishbone_bd_ram_n24670) );
  INV_X1 U31188 ( .A(n62870), .ZN(n26718) );
  INV_X1 U31189 ( .A(n26718), .ZN(p_wishbone_bd_ram_n24669) );
  INV_X1 U31190 ( .A(n62869), .ZN(n26720) );
  INV_X1 U31191 ( .A(n26720), .ZN(p_wishbone_bd_ram_n24668) );
  INV_X1 U31192 ( .A(n62868), .ZN(n26722) );
  INV_X1 U31193 ( .A(n26722), .ZN(p_wishbone_bd_ram_n24667) );
  INV_X1 U31194 ( .A(n62867), .ZN(n26724) );
  INV_X1 U31195 ( .A(n26724), .ZN(p_wishbone_bd_ram_n24666) );
  INV_X1 U31196 ( .A(n62866), .ZN(n26726) );
  INV_X1 U31197 ( .A(n26726), .ZN(p_wishbone_bd_ram_n24665) );
  INV_X1 U31198 ( .A(n62865), .ZN(n26728) );
  INV_X1 U31199 ( .A(n26728), .ZN(p_wishbone_bd_ram_n24664) );
  INV_X1 U31200 ( .A(n62864), .ZN(n26730) );
  INV_X1 U31201 ( .A(n26730), .ZN(p_wishbone_bd_ram_n24663) );
  INV_X1 U31202 ( .A(n62863), .ZN(n26732) );
  INV_X1 U31203 ( .A(n26732), .ZN(p_wishbone_bd_ram_n24662) );
  INV_X1 U31204 ( .A(n62862), .ZN(n26734) );
  INV_X1 U31205 ( .A(n26734), .ZN(p_wishbone_bd_ram_n24661) );
  INV_X1 U31206 ( .A(n62861), .ZN(n26736) );
  INV_X1 U31207 ( .A(n26736), .ZN(p_wishbone_bd_ram_n24660) );
  INV_X1 U31208 ( .A(n62860), .ZN(n26738) );
  INV_X1 U31209 ( .A(n26738), .ZN(p_wishbone_bd_ram_n24659) );
  INV_X1 U31210 ( .A(n62859), .ZN(n26740) );
  INV_X1 U31211 ( .A(n26740), .ZN(p_wishbone_bd_ram_n24658) );
  INV_X1 U31212 ( .A(n62858), .ZN(n26742) );
  INV_X1 U31213 ( .A(n26742), .ZN(p_wishbone_bd_ram_n24657) );
  INV_X1 U31214 ( .A(n62857), .ZN(n26744) );
  INV_X1 U31215 ( .A(n26744), .ZN(p_wishbone_bd_ram_n24656) );
  INV_X1 U31216 ( .A(n62856), .ZN(n26746) );
  INV_X1 U31217 ( .A(n26746), .ZN(p_wishbone_bd_ram_n24655) );
  INV_X1 U31218 ( .A(n62855), .ZN(n26748) );
  INV_X1 U31219 ( .A(n26748), .ZN(p_wishbone_bd_ram_n24654) );
  INV_X1 U31220 ( .A(n62854), .ZN(n26750) );
  INV_X1 U31221 ( .A(n26750), .ZN(p_wishbone_bd_ram_n24653) );
  INV_X1 U31222 ( .A(n62853), .ZN(n26752) );
  INV_X1 U31223 ( .A(n26752), .ZN(p_wishbone_bd_ram_n24652) );
  INV_X1 U31224 ( .A(n62852), .ZN(n26754) );
  INV_X1 U31225 ( .A(n26754), .ZN(p_wishbone_bd_ram_n24651) );
  INV_X1 U31226 ( .A(n62851), .ZN(n26756) );
  INV_X1 U31227 ( .A(n26756), .ZN(p_wishbone_bd_ram_n24650) );
  INV_X1 U31228 ( .A(n62850), .ZN(n26758) );
  INV_X1 U31229 ( .A(n26758), .ZN(p_wishbone_bd_ram_n24649) );
  INV_X1 U31230 ( .A(n62849), .ZN(n26760) );
  INV_X1 U31231 ( .A(n26760), .ZN(p_wishbone_bd_ram_n24648) );
  INV_X1 U31232 ( .A(n62848), .ZN(n26762) );
  INV_X1 U31233 ( .A(n26762), .ZN(p_wishbone_bd_ram_n24647) );
  INV_X1 U31234 ( .A(n62847), .ZN(n26764) );
  INV_X1 U31235 ( .A(n26764), .ZN(p_wishbone_bd_ram_n24646) );
  INV_X1 U31236 ( .A(n62846), .ZN(n26766) );
  INV_X1 U31237 ( .A(n26766), .ZN(p_wishbone_bd_ram_n24645) );
  INV_X1 U31238 ( .A(n62845), .ZN(n26768) );
  INV_X1 U31239 ( .A(n26768), .ZN(p_wishbone_bd_ram_n24644) );
  INV_X1 U31240 ( .A(n62844), .ZN(n26770) );
  INV_X1 U31241 ( .A(n26770), .ZN(p_wishbone_bd_ram_n24643) );
  INV_X1 U31242 ( .A(n62843), .ZN(n26772) );
  INV_X1 U31243 ( .A(n26772), .ZN(p_wishbone_bd_ram_n24642) );
  INV_X1 U31244 ( .A(n62842), .ZN(n26774) );
  INV_X1 U31245 ( .A(n26774), .ZN(p_wishbone_bd_ram_n24641) );
  INV_X1 U31246 ( .A(n62841), .ZN(n26776) );
  INV_X1 U31247 ( .A(n26776), .ZN(p_wishbone_bd_ram_n24640) );
  INV_X1 U31248 ( .A(n62840), .ZN(n26778) );
  INV_X1 U31249 ( .A(n26778), .ZN(p_wishbone_bd_ram_n24639) );
  INV_X1 U31250 ( .A(n62839), .ZN(n26780) );
  INV_X1 U31251 ( .A(n26780), .ZN(p_wishbone_bd_ram_n24638) );
  INV_X1 U31252 ( .A(n62838), .ZN(n26782) );
  INV_X1 U31253 ( .A(n26782), .ZN(p_wishbone_bd_ram_n24637) );
  INV_X1 U31254 ( .A(n62837), .ZN(n26784) );
  INV_X1 U31255 ( .A(n26784), .ZN(p_wishbone_bd_ram_n24636) );
  INV_X1 U31256 ( .A(n62836), .ZN(n26786) );
  INV_X1 U31257 ( .A(n26786), .ZN(p_wishbone_bd_ram_n24635) );
  INV_X1 U31258 ( .A(n62835), .ZN(n26788) );
  INV_X1 U31259 ( .A(n26788), .ZN(p_wishbone_bd_ram_n24634) );
  INV_X1 U31260 ( .A(n62834), .ZN(n26790) );
  INV_X1 U31261 ( .A(n26790), .ZN(p_wishbone_bd_ram_n24633) );
  INV_X1 U31262 ( .A(n62833), .ZN(n26792) );
  INV_X1 U31263 ( .A(n26792), .ZN(p_wishbone_bd_ram_n24632) );
  INV_X1 U31264 ( .A(n62832), .ZN(n26794) );
  INV_X1 U31265 ( .A(n26794), .ZN(p_wishbone_bd_ram_n24631) );
  INV_X1 U31266 ( .A(n62831), .ZN(n26796) );
  INV_X1 U31267 ( .A(n26796), .ZN(p_wishbone_bd_ram_n24630) );
  INV_X1 U31268 ( .A(n62830), .ZN(n26798) );
  INV_X1 U31269 ( .A(n26798), .ZN(p_wishbone_bd_ram_n24629) );
  INV_X1 U31270 ( .A(n62829), .ZN(n26800) );
  INV_X1 U31271 ( .A(n26800), .ZN(p_wishbone_bd_ram_n24628) );
  INV_X1 U31272 ( .A(n62828), .ZN(n26802) );
  INV_X1 U31273 ( .A(n26802), .ZN(p_wishbone_bd_ram_n24627) );
  INV_X1 U31274 ( .A(n62827), .ZN(n26804) );
  INV_X1 U31275 ( .A(n26804), .ZN(p_wishbone_bd_ram_n24626) );
  INV_X1 U31276 ( .A(n62826), .ZN(n26806) );
  INV_X1 U31277 ( .A(n26806), .ZN(p_wishbone_bd_ram_n24625) );
  INV_X1 U31278 ( .A(n62825), .ZN(n26808) );
  INV_X1 U31279 ( .A(n26808), .ZN(p_wishbone_bd_ram_n24624) );
  INV_X1 U31280 ( .A(n62824), .ZN(n26810) );
  INV_X1 U31281 ( .A(n26810), .ZN(p_wishbone_bd_ram_n24623) );
  INV_X1 U31282 ( .A(n62823), .ZN(n26812) );
  INV_X1 U31283 ( .A(n26812), .ZN(p_wishbone_bd_ram_n24622) );
  INV_X1 U31284 ( .A(n62822), .ZN(n26814) );
  INV_X1 U31285 ( .A(n26814), .ZN(p_wishbone_bd_ram_n24621) );
  INV_X1 U31286 ( .A(n62821), .ZN(n26816) );
  INV_X1 U31287 ( .A(n26816), .ZN(p_wishbone_bd_ram_n24620) );
  INV_X1 U31288 ( .A(n62820), .ZN(n26818) );
  INV_X1 U31289 ( .A(n26818), .ZN(p_wishbone_bd_ram_n24619) );
  INV_X1 U31290 ( .A(n62819), .ZN(n26820) );
  INV_X1 U31291 ( .A(n26820), .ZN(p_wishbone_bd_ram_n24618) );
  INV_X1 U31292 ( .A(n62818), .ZN(n26822) );
  INV_X1 U31293 ( .A(n26822), .ZN(p_wishbone_bd_ram_n24617) );
  INV_X1 U31294 ( .A(n62817), .ZN(n26824) );
  INV_X1 U31295 ( .A(n26824), .ZN(p_wishbone_bd_ram_n24616) );
  INV_X1 U31296 ( .A(n62816), .ZN(n26826) );
  INV_X1 U31297 ( .A(n26826), .ZN(p_wishbone_bd_ram_n24615) );
  INV_X1 U31298 ( .A(n62815), .ZN(n26828) );
  INV_X1 U31299 ( .A(n26828), .ZN(p_wishbone_bd_ram_n24614) );
  INV_X1 U31300 ( .A(n62814), .ZN(n26830) );
  INV_X1 U31301 ( .A(n26830), .ZN(p_wishbone_bd_ram_n24613) );
  INV_X1 U31302 ( .A(n62813), .ZN(n26832) );
  INV_X1 U31303 ( .A(n26832), .ZN(p_wishbone_bd_ram_n24612) );
  INV_X1 U31304 ( .A(n62812), .ZN(n26834) );
  INV_X1 U31305 ( .A(n26834), .ZN(p_wishbone_bd_ram_n24611) );
  INV_X1 U31306 ( .A(n62811), .ZN(n26836) );
  INV_X1 U31307 ( .A(n26836), .ZN(p_wishbone_bd_ram_n24610) );
  INV_X1 U31308 ( .A(n62810), .ZN(n26838) );
  INV_X1 U31309 ( .A(n26838), .ZN(p_wishbone_bd_ram_n24609) );
  INV_X1 U31310 ( .A(n62809), .ZN(n26840) );
  INV_X1 U31311 ( .A(n26840), .ZN(p_wishbone_bd_ram_n24607) );
  INV_X1 U31312 ( .A(n62808), .ZN(n26842) );
  INV_X1 U31313 ( .A(n26842), .ZN(p_wishbone_bd_ram_n24605) );
  INV_X1 U31314 ( .A(n62807), .ZN(n26844) );
  INV_X1 U31315 ( .A(n26844), .ZN(p_wishbone_bd_ram_n24604) );
  INV_X1 U31316 ( .A(n62806), .ZN(n26846) );
  INV_X1 U31317 ( .A(n26846), .ZN(p_wishbone_bd_ram_n24602) );
  INV_X1 U31318 ( .A(n62805), .ZN(n26848) );
  INV_X1 U31319 ( .A(n26848), .ZN(p_wishbone_bd_ram_n24600) );
  INV_X1 U31320 ( .A(n62804), .ZN(n26850) );
  INV_X1 U31321 ( .A(n26850), .ZN(p_wishbone_bd_ram_n24599) );
  INV_X1 U31322 ( .A(n62803), .ZN(n26852) );
  INV_X1 U31323 ( .A(n26852), .ZN(p_wishbone_bd_ram_n24598) );
  INV_X1 U31324 ( .A(n62802), .ZN(n26854) );
  INV_X1 U31325 ( .A(n26854), .ZN(p_wishbone_bd_ram_n24597) );
  INV_X1 U31326 ( .A(n62801), .ZN(n26856) );
  INV_X1 U31327 ( .A(n26856), .ZN(p_wishbone_bd_ram_n24596) );
  INV_X1 U31328 ( .A(n62800), .ZN(n26858) );
  INV_X1 U31329 ( .A(n26858), .ZN(p_wishbone_bd_ram_n24595) );
  INV_X1 U31330 ( .A(n62799), .ZN(n26860) );
  INV_X1 U31331 ( .A(n26860), .ZN(p_wishbone_bd_ram_n24594) );
  INV_X1 U31332 ( .A(n62798), .ZN(n26862) );
  INV_X1 U31333 ( .A(n26862), .ZN(p_wishbone_bd_ram_n24593) );
  INV_X1 U31334 ( .A(n62797), .ZN(n26864) );
  INV_X1 U31335 ( .A(n26864), .ZN(p_wishbone_bd_ram_n24592) );
  INV_X1 U31336 ( .A(n62796), .ZN(n26866) );
  INV_X1 U31337 ( .A(n26866), .ZN(p_wishbone_bd_ram_n24591) );
  INV_X1 U31338 ( .A(n62795), .ZN(n26868) );
  INV_X1 U31339 ( .A(n26868), .ZN(p_wishbone_bd_ram_n24590) );
  INV_X1 U31340 ( .A(n62794), .ZN(n26870) );
  INV_X1 U31341 ( .A(n26870), .ZN(p_wishbone_bd_ram_n24589) );
  INV_X1 U31342 ( .A(n62793), .ZN(n26872) );
  INV_X1 U31343 ( .A(n26872), .ZN(p_wishbone_bd_ram_n24588) );
  INV_X1 U31344 ( .A(n62792), .ZN(n26874) );
  INV_X1 U31345 ( .A(n26874), .ZN(p_wishbone_bd_ram_n24587) );
  INV_X1 U31346 ( .A(n62791), .ZN(n26876) );
  INV_X1 U31347 ( .A(n26876), .ZN(p_wishbone_bd_ram_n24586) );
  INV_X1 U31348 ( .A(n62790), .ZN(n26878) );
  INV_X1 U31349 ( .A(n26878), .ZN(p_wishbone_bd_ram_n24585) );
  INV_X1 U31350 ( .A(n62789), .ZN(n26880) );
  INV_X1 U31351 ( .A(n26880), .ZN(p_wishbone_bd_ram_n24583) );
  INV_X1 U31352 ( .A(n62788), .ZN(n26882) );
  INV_X1 U31353 ( .A(n26882), .ZN(p_wishbone_bd_ram_n24581) );
  INV_X1 U31354 ( .A(n62787), .ZN(n26884) );
  INV_X1 U31355 ( .A(n26884), .ZN(p_wishbone_bd_ram_n24580) );
  INV_X1 U31356 ( .A(n62786), .ZN(n26886) );
  INV_X1 U31357 ( .A(n26886), .ZN(p_wishbone_bd_ram_n24578) );
  INV_X1 U31358 ( .A(n62785), .ZN(n26888) );
  INV_X1 U31359 ( .A(n26888), .ZN(p_wishbone_bd_ram_n24576) );
  INV_X1 U31360 ( .A(n62784), .ZN(n26890) );
  INV_X1 U31361 ( .A(n26890), .ZN(p_wishbone_bd_ram_n24575) );
  INV_X1 U31362 ( .A(n62783), .ZN(n26892) );
  INV_X1 U31363 ( .A(n26892), .ZN(p_wishbone_bd_ram_n24574) );
  INV_X1 U31364 ( .A(n62782), .ZN(n26894) );
  INV_X1 U31365 ( .A(n26894), .ZN(p_wishbone_bd_ram_n24573) );
  INV_X1 U31366 ( .A(n62781), .ZN(n26896) );
  INV_X1 U31367 ( .A(n26896), .ZN(p_wishbone_bd_ram_n24572) );
  INV_X1 U31368 ( .A(n62780), .ZN(n26898) );
  INV_X1 U31369 ( .A(n26898), .ZN(p_wishbone_bd_ram_n24571) );
  INV_X1 U31370 ( .A(n62779), .ZN(n26900) );
  INV_X1 U31371 ( .A(n26900), .ZN(p_wishbone_bd_ram_n24570) );
  INV_X1 U31372 ( .A(n62778), .ZN(n26902) );
  INV_X1 U31373 ( .A(n26902), .ZN(p_wishbone_bd_ram_n24569) );
  INV_X1 U31374 ( .A(n62777), .ZN(n26904) );
  INV_X1 U31375 ( .A(n26904), .ZN(p_wishbone_bd_ram_n24568) );
  INV_X1 U31376 ( .A(n62776), .ZN(n26906) );
  INV_X1 U31377 ( .A(n26906), .ZN(p_wishbone_bd_ram_n24567) );
  INV_X1 U31378 ( .A(n62775), .ZN(n26908) );
  INV_X1 U31379 ( .A(n26908), .ZN(p_wishbone_bd_ram_n24566) );
  INV_X1 U31380 ( .A(n62774), .ZN(n26910) );
  INV_X1 U31381 ( .A(n26910), .ZN(p_wishbone_bd_ram_n24565) );
  INV_X1 U31382 ( .A(n62773), .ZN(n26912) );
  INV_X1 U31383 ( .A(n26912), .ZN(p_wishbone_bd_ram_n24564) );
  INV_X1 U31384 ( .A(n62772), .ZN(n26914) );
  INV_X1 U31385 ( .A(n26914), .ZN(p_wishbone_bd_ram_n24563) );
  INV_X1 U31386 ( .A(n62771), .ZN(n26916) );
  INV_X1 U31387 ( .A(n26916), .ZN(p_wishbone_bd_ram_n24562) );
  INV_X1 U31388 ( .A(n62770), .ZN(n26918) );
  INV_X1 U31389 ( .A(n26918), .ZN(p_wishbone_bd_ram_n24561) );
  INV_X1 U31390 ( .A(n62769), .ZN(n26920) );
  INV_X1 U31391 ( .A(n26920), .ZN(p_wishbone_bd_ram_n24560) );
  INV_X1 U31392 ( .A(n62768), .ZN(n26922) );
  INV_X1 U31393 ( .A(n26922), .ZN(p_wishbone_bd_ram_n24559) );
  INV_X1 U31394 ( .A(n62767), .ZN(n26924) );
  INV_X1 U31395 ( .A(n26924), .ZN(p_wishbone_bd_ram_n24558) );
  INV_X1 U31396 ( .A(n62766), .ZN(n26926) );
  INV_X1 U31397 ( .A(n26926), .ZN(p_wishbone_bd_ram_n24557) );
  INV_X1 U31398 ( .A(n62765), .ZN(n26928) );
  INV_X1 U31399 ( .A(n26928), .ZN(p_wishbone_bd_ram_n24556) );
  INV_X1 U31400 ( .A(n62764), .ZN(n26930) );
  INV_X1 U31401 ( .A(n26930), .ZN(p_wishbone_bd_ram_n24555) );
  INV_X1 U31402 ( .A(n62763), .ZN(n26932) );
  INV_X1 U31403 ( .A(n26932), .ZN(p_wishbone_bd_ram_n24554) );
  INV_X1 U31404 ( .A(n62762), .ZN(n26934) );
  INV_X1 U31405 ( .A(n26934), .ZN(p_wishbone_bd_ram_n24553) );
  INV_X1 U31406 ( .A(n62761), .ZN(n26936) );
  INV_X1 U31407 ( .A(n26936), .ZN(p_wishbone_bd_ram_n24552) );
  INV_X1 U31408 ( .A(n62760), .ZN(n26938) );
  INV_X1 U31409 ( .A(n26938), .ZN(p_wishbone_bd_ram_n24551) );
  INV_X1 U31410 ( .A(n62759), .ZN(n26940) );
  INV_X1 U31411 ( .A(n26940), .ZN(p_wishbone_bd_ram_n24550) );
  INV_X1 U31412 ( .A(n62758), .ZN(n26942) );
  INV_X1 U31413 ( .A(n26942), .ZN(p_wishbone_bd_ram_n24549) );
  INV_X1 U31414 ( .A(n62757), .ZN(n26944) );
  INV_X1 U31415 ( .A(n26944), .ZN(p_wishbone_bd_ram_n24548) );
  INV_X1 U31416 ( .A(n62756), .ZN(n26946) );
  INV_X1 U31417 ( .A(n26946), .ZN(p_wishbone_bd_ram_n24547) );
  INV_X1 U31418 ( .A(n62755), .ZN(n26948) );
  INV_X1 U31419 ( .A(n26948), .ZN(p_wishbone_bd_ram_n24546) );
  INV_X1 U31420 ( .A(n62754), .ZN(n26950) );
  INV_X1 U31421 ( .A(n26950), .ZN(p_wishbone_bd_ram_n24545) );
  INV_X1 U31422 ( .A(n62753), .ZN(n26952) );
  INV_X1 U31423 ( .A(n26952), .ZN(p_wishbone_bd_ram_n24544) );
  INV_X1 U31424 ( .A(n62752), .ZN(n26954) );
  INV_X1 U31425 ( .A(n26954), .ZN(p_wishbone_bd_ram_n24543) );
  INV_X1 U31426 ( .A(n62751), .ZN(n26956) );
  INV_X1 U31427 ( .A(n26956), .ZN(p_wishbone_bd_ram_n24542) );
  INV_X1 U31428 ( .A(n62750), .ZN(n26958) );
  INV_X1 U31429 ( .A(n26958), .ZN(p_wishbone_bd_ram_n24541) );
  INV_X1 U31430 ( .A(n62749), .ZN(n26960) );
  INV_X1 U31431 ( .A(n26960), .ZN(p_wishbone_bd_ram_n24540) );
  INV_X1 U31432 ( .A(n62748), .ZN(n26962) );
  INV_X1 U31433 ( .A(n26962), .ZN(p_wishbone_bd_ram_n24539) );
  INV_X1 U31434 ( .A(n62747), .ZN(n26964) );
  INV_X1 U31435 ( .A(n26964), .ZN(p_wishbone_bd_ram_n24538) );
  INV_X1 U31436 ( .A(n62746), .ZN(n26966) );
  INV_X1 U31437 ( .A(n26966), .ZN(p_wishbone_bd_ram_n24537) );
  INV_X1 U31438 ( .A(n62745), .ZN(n26968) );
  INV_X1 U31439 ( .A(n26968), .ZN(p_wishbone_bd_ram_n24536) );
  INV_X1 U31440 ( .A(n62744), .ZN(n26970) );
  INV_X1 U31441 ( .A(n26970), .ZN(p_wishbone_bd_ram_n24535) );
  INV_X1 U31442 ( .A(n62743), .ZN(n26972) );
  INV_X1 U31443 ( .A(n26972), .ZN(p_wishbone_bd_ram_n24534) );
  INV_X1 U31444 ( .A(n62742), .ZN(n26974) );
  INV_X1 U31445 ( .A(n26974), .ZN(p_wishbone_bd_ram_n24533) );
  INV_X1 U31446 ( .A(n62741), .ZN(n26976) );
  INV_X1 U31447 ( .A(n26976), .ZN(p_wishbone_bd_ram_n24532) );
  INV_X1 U31448 ( .A(n62740), .ZN(n26978) );
  INV_X1 U31449 ( .A(n26978), .ZN(p_wishbone_bd_ram_n24531) );
  INV_X1 U31450 ( .A(n62739), .ZN(n26980) );
  INV_X1 U31451 ( .A(n26980), .ZN(p_wishbone_bd_ram_n24530) );
  INV_X1 U31452 ( .A(n62738), .ZN(n26982) );
  INV_X1 U31453 ( .A(n26982), .ZN(p_wishbone_bd_ram_n24529) );
  INV_X1 U31454 ( .A(n62737), .ZN(n26984) );
  INV_X1 U31455 ( .A(n26984), .ZN(p_wishbone_bd_ram_n24527) );
  INV_X1 U31456 ( .A(n62736), .ZN(n26986) );
  INV_X1 U31457 ( .A(n26986), .ZN(p_wishbone_bd_ram_n24525) );
  INV_X1 U31458 ( .A(n62735), .ZN(n26988) );
  INV_X1 U31459 ( .A(n26988), .ZN(p_wishbone_bd_ram_n24524) );
  INV_X1 U31460 ( .A(n62734), .ZN(n26990) );
  INV_X1 U31461 ( .A(n26990), .ZN(p_wishbone_bd_ram_n24522) );
  INV_X1 U31462 ( .A(n62733), .ZN(n26992) );
  INV_X1 U31463 ( .A(n26992), .ZN(p_wishbone_bd_ram_n24519) );
  INV_X1 U31464 ( .A(n62732), .ZN(n26994) );
  INV_X1 U31465 ( .A(n26994), .ZN(p_wishbone_bd_ram_n24517) );
  INV_X1 U31466 ( .A(n62731), .ZN(n26996) );
  INV_X1 U31467 ( .A(n26996), .ZN(p_wishbone_bd_ram_n24516) );
  INV_X1 U31468 ( .A(n62730), .ZN(n26998) );
  INV_X1 U31469 ( .A(n26998), .ZN(p_wishbone_bd_ram_n24514) );
  INV_X1 U31470 ( .A(n62729), .ZN(n27000) );
  INV_X1 U31471 ( .A(n27000), .ZN(p_wishbone_bd_ram_n24512) );
  INV_X1 U31472 ( .A(n62728), .ZN(n27002) );
  INV_X1 U31473 ( .A(n27002), .ZN(p_wishbone_bd_ram_n24511) );
  INV_X1 U31474 ( .A(n62727), .ZN(n27004) );
  INV_X1 U31475 ( .A(n27004), .ZN(p_wishbone_bd_ram_n24510) );
  INV_X1 U31476 ( .A(n62726), .ZN(n27006) );
  INV_X1 U31477 ( .A(n27006), .ZN(p_wishbone_bd_ram_n24509) );
  INV_X1 U31478 ( .A(n62725), .ZN(n27008) );
  INV_X1 U31479 ( .A(n27008), .ZN(p_wishbone_bd_ram_n24508) );
  INV_X1 U31480 ( .A(n62724), .ZN(n27010) );
  INV_X1 U31481 ( .A(n27010), .ZN(p_wishbone_bd_ram_n24507) );
  INV_X1 U31482 ( .A(n62723), .ZN(n27012) );
  INV_X1 U31483 ( .A(n27012), .ZN(p_wishbone_bd_ram_n24506) );
  INV_X1 U31484 ( .A(n62722), .ZN(n27014) );
  INV_X1 U31485 ( .A(n27014), .ZN(p_wishbone_bd_ram_n24505) );
  INV_X1 U31486 ( .A(n62721), .ZN(n27016) );
  INV_X1 U31487 ( .A(n27016), .ZN(p_wishbone_bd_ram_n24504) );
  INV_X1 U31488 ( .A(n62720), .ZN(n27018) );
  INV_X1 U31489 ( .A(n27018), .ZN(p_wishbone_bd_ram_n24503) );
  INV_X1 U31490 ( .A(n62719), .ZN(n27020) );
  INV_X1 U31491 ( .A(n27020), .ZN(p_wishbone_bd_ram_n24502) );
  INV_X1 U31492 ( .A(n62718), .ZN(n27022) );
  INV_X1 U31493 ( .A(n27022), .ZN(p_wishbone_bd_ram_n24501) );
  INV_X1 U31494 ( .A(n62717), .ZN(n27024) );
  INV_X1 U31495 ( .A(n27024), .ZN(p_wishbone_bd_ram_n24500) );
  INV_X1 U31496 ( .A(n62716), .ZN(n27026) );
  INV_X1 U31497 ( .A(n27026), .ZN(p_wishbone_bd_ram_n24499) );
  INV_X1 U31498 ( .A(n62715), .ZN(n27028) );
  INV_X1 U31499 ( .A(n27028), .ZN(p_wishbone_bd_ram_n24498) );
  INV_X1 U31500 ( .A(n62714), .ZN(n27030) );
  INV_X1 U31501 ( .A(n27030), .ZN(p_wishbone_bd_ram_n24497) );
  INV_X1 U31502 ( .A(n62713), .ZN(n27032) );
  INV_X1 U31503 ( .A(n27032), .ZN(p_wishbone_bd_ram_n24496) );
  INV_X1 U31504 ( .A(n62712), .ZN(n27034) );
  INV_X1 U31505 ( .A(n27034), .ZN(p_wishbone_bd_ram_n24495) );
  INV_X1 U31506 ( .A(n62711), .ZN(n27036) );
  INV_X1 U31507 ( .A(n27036), .ZN(p_wishbone_bd_ram_n24494) );
  INV_X1 U31508 ( .A(n62710), .ZN(n27038) );
  INV_X1 U31509 ( .A(n27038), .ZN(p_wishbone_bd_ram_n24493) );
  INV_X1 U31510 ( .A(n62709), .ZN(n27040) );
  INV_X1 U31511 ( .A(n27040), .ZN(p_wishbone_bd_ram_n24492) );
  INV_X1 U31512 ( .A(n62708), .ZN(n27042) );
  INV_X1 U31513 ( .A(n27042), .ZN(p_wishbone_bd_ram_n24491) );
  INV_X1 U31514 ( .A(n62707), .ZN(n27044) );
  INV_X1 U31515 ( .A(n27044), .ZN(p_wishbone_bd_ram_n24490) );
  INV_X1 U31516 ( .A(n62706), .ZN(n27046) );
  INV_X1 U31517 ( .A(n27046), .ZN(p_wishbone_bd_ram_n24489) );
  INV_X1 U31518 ( .A(n62705), .ZN(n27048) );
  INV_X1 U31519 ( .A(n27048), .ZN(p_wishbone_bd_ram_n24488) );
  INV_X1 U31520 ( .A(n62704), .ZN(n27050) );
  INV_X1 U31521 ( .A(n27050), .ZN(p_wishbone_bd_ram_n24487) );
  INV_X1 U31522 ( .A(n62703), .ZN(n27052) );
  INV_X1 U31523 ( .A(n27052), .ZN(p_wishbone_bd_ram_n24486) );
  INV_X1 U31524 ( .A(n62702), .ZN(n27054) );
  INV_X1 U31525 ( .A(n27054), .ZN(p_wishbone_bd_ram_n24485) );
  INV_X1 U31526 ( .A(n62701), .ZN(n27056) );
  INV_X1 U31527 ( .A(n27056), .ZN(p_wishbone_bd_ram_n24484) );
  INV_X1 U31528 ( .A(n62700), .ZN(n27058) );
  INV_X1 U31529 ( .A(n27058), .ZN(p_wishbone_bd_ram_n24483) );
  INV_X1 U31530 ( .A(n62699), .ZN(n27060) );
  INV_X1 U31531 ( .A(n27060), .ZN(p_wishbone_bd_ram_n24482) );
  INV_X1 U31532 ( .A(n62698), .ZN(n27062) );
  INV_X1 U31533 ( .A(n27062), .ZN(p_wishbone_bd_ram_n24481) );
  INV_X1 U31534 ( .A(n62697), .ZN(n27064) );
  INV_X1 U31535 ( .A(n27064), .ZN(p_wishbone_bd_ram_n24480) );
  INV_X1 U31536 ( .A(n62696), .ZN(n27066) );
  INV_X1 U31537 ( .A(n27066), .ZN(p_wishbone_bd_ram_n24479) );
  INV_X1 U31538 ( .A(n62695), .ZN(n27068) );
  INV_X1 U31539 ( .A(n27068), .ZN(p_wishbone_bd_ram_n24478) );
  INV_X1 U31540 ( .A(n62694), .ZN(n27070) );
  INV_X1 U31541 ( .A(n27070), .ZN(p_wishbone_bd_ram_n24477) );
  INV_X1 U31542 ( .A(n62693), .ZN(n27072) );
  INV_X1 U31543 ( .A(n27072), .ZN(p_wishbone_bd_ram_n24476) );
  INV_X1 U31544 ( .A(n62692), .ZN(n27074) );
  INV_X1 U31545 ( .A(n27074), .ZN(p_wishbone_bd_ram_n24475) );
  INV_X1 U31546 ( .A(n62691), .ZN(n27076) );
  INV_X1 U31547 ( .A(n27076), .ZN(p_wishbone_bd_ram_n24474) );
  INV_X1 U31548 ( .A(n62690), .ZN(n27078) );
  INV_X1 U31549 ( .A(n27078), .ZN(p_wishbone_bd_ram_n24473) );
  INV_X1 U31550 ( .A(n62689), .ZN(n27080) );
  INV_X1 U31551 ( .A(n27080), .ZN(p_wishbone_bd_ram_n24472) );
  INV_X1 U31552 ( .A(n62688), .ZN(n27082) );
  INV_X1 U31553 ( .A(n27082), .ZN(p_wishbone_bd_ram_n24471) );
  INV_X1 U31554 ( .A(n62687), .ZN(n27084) );
  INV_X1 U31555 ( .A(n27084), .ZN(p_wishbone_bd_ram_n24470) );
  INV_X1 U31556 ( .A(n62686), .ZN(n27086) );
  INV_X1 U31557 ( .A(n27086), .ZN(p_wishbone_bd_ram_n24469) );
  INV_X1 U31558 ( .A(n62685), .ZN(n27088) );
  INV_X1 U31559 ( .A(n27088), .ZN(p_wishbone_bd_ram_n24468) );
  INV_X1 U31560 ( .A(n62684), .ZN(n27090) );
  INV_X1 U31561 ( .A(n27090), .ZN(p_wishbone_bd_ram_n24467) );
  INV_X1 U31562 ( .A(n62683), .ZN(n27092) );
  INV_X1 U31563 ( .A(n27092), .ZN(p_wishbone_bd_ram_n24466) );
  INV_X1 U31564 ( .A(n62682), .ZN(n27094) );
  INV_X1 U31565 ( .A(n27094), .ZN(p_wishbone_bd_ram_n24465) );
  INV_X1 U31566 ( .A(n62681), .ZN(n27096) );
  INV_X1 U31567 ( .A(n27096), .ZN(p_wishbone_bd_ram_n24464) );
  INV_X1 U31568 ( .A(n62680), .ZN(n27098) );
  INV_X1 U31569 ( .A(n27098), .ZN(p_wishbone_bd_ram_n24463) );
  INV_X1 U31570 ( .A(n62679), .ZN(n27100) );
  INV_X1 U31571 ( .A(n27100), .ZN(p_wishbone_bd_ram_n24462) );
  INV_X1 U31572 ( .A(n62678), .ZN(n27102) );
  INV_X1 U31573 ( .A(n27102), .ZN(p_wishbone_bd_ram_n24461) );
  INV_X1 U31574 ( .A(n62677), .ZN(n27104) );
  INV_X1 U31575 ( .A(n27104), .ZN(p_wishbone_bd_ram_n24460) );
  INV_X1 U31576 ( .A(n62676), .ZN(n27106) );
  INV_X1 U31577 ( .A(n27106), .ZN(p_wishbone_bd_ram_n24459) );
  INV_X1 U31578 ( .A(n62675), .ZN(n27108) );
  INV_X1 U31579 ( .A(n27108), .ZN(p_wishbone_bd_ram_n24458) );
  INV_X1 U31580 ( .A(n62674), .ZN(n27110) );
  INV_X1 U31581 ( .A(n27110), .ZN(p_wishbone_bd_ram_n24457) );
  INV_X1 U31582 ( .A(n62673), .ZN(n27112) );
  INV_X1 U31583 ( .A(n27112), .ZN(p_wishbone_bd_ram_n24456) );
  INV_X1 U31584 ( .A(n62672), .ZN(n27114) );
  INV_X1 U31585 ( .A(n27114), .ZN(p_wishbone_bd_ram_n24455) );
  INV_X1 U31586 ( .A(n62671), .ZN(n27116) );
  INV_X1 U31587 ( .A(n27116), .ZN(p_wishbone_bd_ram_n24454) );
  INV_X1 U31588 ( .A(n62670), .ZN(n27118) );
  INV_X1 U31589 ( .A(n27118), .ZN(p_wishbone_bd_ram_n24453) );
  INV_X1 U31590 ( .A(n62669), .ZN(n27120) );
  INV_X1 U31591 ( .A(n27120), .ZN(p_wishbone_bd_ram_n24452) );
  INV_X1 U31592 ( .A(n62668), .ZN(n27122) );
  INV_X1 U31593 ( .A(n27122), .ZN(p_wishbone_bd_ram_n24451) );
  INV_X1 U31594 ( .A(n62667), .ZN(n27124) );
  INV_X1 U31595 ( .A(n27124), .ZN(p_wishbone_bd_ram_n24450) );
  INV_X1 U31596 ( .A(n62666), .ZN(n27126) );
  INV_X1 U31597 ( .A(n27126), .ZN(p_wishbone_bd_ram_n24449) );
  INV_X1 U31598 ( .A(n62665), .ZN(n27128) );
  INV_X1 U31599 ( .A(n27128), .ZN(p_wishbone_bd_ram_n24448) );
  INV_X1 U31600 ( .A(n62664), .ZN(n27130) );
  INV_X1 U31601 ( .A(n27130), .ZN(p_wishbone_bd_ram_n24447) );
  INV_X1 U31602 ( .A(n62663), .ZN(n27132) );
  INV_X1 U31603 ( .A(n27132), .ZN(p_wishbone_bd_ram_n24446) );
  INV_X1 U31604 ( .A(n62662), .ZN(n27134) );
  INV_X1 U31605 ( .A(n27134), .ZN(p_wishbone_bd_ram_n24445) );
  INV_X1 U31606 ( .A(n62661), .ZN(n27136) );
  INV_X1 U31607 ( .A(n27136), .ZN(p_wishbone_bd_ram_n24444) );
  INV_X1 U31608 ( .A(n62660), .ZN(n27138) );
  INV_X1 U31609 ( .A(n27138), .ZN(p_wishbone_bd_ram_n24443) );
  INV_X1 U31610 ( .A(n62659), .ZN(n27140) );
  INV_X1 U31611 ( .A(n27140), .ZN(p_wishbone_bd_ram_n24442) );
  INV_X1 U31612 ( .A(n62658), .ZN(n27142) );
  INV_X1 U31613 ( .A(n27142), .ZN(p_wishbone_bd_ram_n24441) );
  INV_X1 U31614 ( .A(n62657), .ZN(n27144) );
  INV_X1 U31615 ( .A(n27144), .ZN(p_wishbone_bd_ram_n24440) );
  INV_X1 U31616 ( .A(n62656), .ZN(n27146) );
  INV_X1 U31617 ( .A(n27146), .ZN(p_wishbone_bd_ram_n24439) );
  INV_X1 U31618 ( .A(n62655), .ZN(n27148) );
  INV_X1 U31619 ( .A(n27148), .ZN(p_wishbone_bd_ram_n24438) );
  INV_X1 U31620 ( .A(n62654), .ZN(n27150) );
  INV_X1 U31621 ( .A(n27150), .ZN(p_wishbone_bd_ram_n24437) );
  INV_X1 U31622 ( .A(n62653), .ZN(n27152) );
  INV_X1 U31623 ( .A(n27152), .ZN(p_wishbone_bd_ram_n24436) );
  INV_X1 U31624 ( .A(n62652), .ZN(n27154) );
  INV_X1 U31625 ( .A(n27154), .ZN(p_wishbone_bd_ram_n24435) );
  INV_X1 U31626 ( .A(n62651), .ZN(n27156) );
  INV_X1 U31627 ( .A(n27156), .ZN(p_wishbone_bd_ram_n24434) );
  INV_X1 U31628 ( .A(n62650), .ZN(n27158) );
  INV_X1 U31629 ( .A(n27158), .ZN(p_wishbone_bd_ram_n24433) );
  INV_X1 U31630 ( .A(n62649), .ZN(n27160) );
  INV_X1 U31631 ( .A(n27160), .ZN(p_wishbone_bd_ram_n24432) );
  INV_X1 U31632 ( .A(n62648), .ZN(n27162) );
  INV_X1 U31633 ( .A(n27162), .ZN(p_wishbone_bd_ram_n24431) );
  INV_X1 U31634 ( .A(n62647), .ZN(n27164) );
  INV_X1 U31635 ( .A(n27164), .ZN(p_wishbone_bd_ram_n24430) );
  INV_X1 U31636 ( .A(n62646), .ZN(n27166) );
  INV_X1 U31637 ( .A(n27166), .ZN(p_wishbone_bd_ram_n24429) );
  INV_X1 U31638 ( .A(n62645), .ZN(n27168) );
  INV_X1 U31639 ( .A(n27168), .ZN(p_wishbone_bd_ram_n24428) );
  INV_X1 U31640 ( .A(n62644), .ZN(n27170) );
  INV_X1 U31641 ( .A(n27170), .ZN(p_wishbone_bd_ram_n24427) );
  INV_X1 U31642 ( .A(n62643), .ZN(n27172) );
  INV_X1 U31643 ( .A(n27172), .ZN(p_wishbone_bd_ram_n24426) );
  INV_X1 U31644 ( .A(n62642), .ZN(n27174) );
  INV_X1 U31645 ( .A(n27174), .ZN(p_wishbone_bd_ram_n24425) );
  INV_X1 U31646 ( .A(n62641), .ZN(n27176) );
  INV_X1 U31647 ( .A(n27176), .ZN(p_wishbone_bd_ram_n24424) );
  INV_X1 U31648 ( .A(n62640), .ZN(n27178) );
  INV_X1 U31649 ( .A(n27178), .ZN(p_wishbone_bd_ram_n24423) );
  INV_X1 U31650 ( .A(n62639), .ZN(n27180) );
  INV_X1 U31651 ( .A(n27180), .ZN(p_wishbone_bd_ram_n24422) );
  INV_X1 U31652 ( .A(n62638), .ZN(n27182) );
  INV_X1 U31653 ( .A(n27182), .ZN(p_wishbone_bd_ram_n24421) );
  INV_X1 U31654 ( .A(n62637), .ZN(n27184) );
  INV_X1 U31655 ( .A(n27184), .ZN(p_wishbone_bd_ram_n24420) );
  INV_X1 U31656 ( .A(n62636), .ZN(n27186) );
  INV_X1 U31657 ( .A(n27186), .ZN(p_wishbone_bd_ram_n24419) );
  INV_X1 U31658 ( .A(n62635), .ZN(n27188) );
  INV_X1 U31659 ( .A(n27188), .ZN(p_wishbone_bd_ram_n24418) );
  INV_X1 U31660 ( .A(n62634), .ZN(n27190) );
  INV_X1 U31661 ( .A(n27190), .ZN(p_wishbone_bd_ram_n24417) );
  INV_X1 U31662 ( .A(n62633), .ZN(n27192) );
  INV_X1 U31663 ( .A(n27192), .ZN(p_wishbone_bd_ram_n24416) );
  INV_X1 U31664 ( .A(n62632), .ZN(n27194) );
  INV_X1 U31665 ( .A(n27194), .ZN(p_wishbone_bd_ram_n24415) );
  INV_X1 U31666 ( .A(n62631), .ZN(n27196) );
  INV_X1 U31667 ( .A(n27196), .ZN(p_wishbone_bd_ram_n24414) );
  INV_X1 U31668 ( .A(n62630), .ZN(n27198) );
  INV_X1 U31669 ( .A(n27198), .ZN(p_wishbone_bd_ram_n24413) );
  INV_X1 U31670 ( .A(n62629), .ZN(n27200) );
  INV_X1 U31671 ( .A(n27200), .ZN(p_wishbone_bd_ram_n24412) );
  INV_X1 U31672 ( .A(n62628), .ZN(n27202) );
  INV_X1 U31673 ( .A(n27202), .ZN(p_wishbone_bd_ram_n24411) );
  INV_X1 U31674 ( .A(n62627), .ZN(n27204) );
  INV_X1 U31675 ( .A(n27204), .ZN(p_wishbone_bd_ram_n24410) );
  INV_X1 U31676 ( .A(n62626), .ZN(n27206) );
  INV_X1 U31677 ( .A(n27206), .ZN(p_wishbone_bd_ram_n24409) );
  INV_X1 U31678 ( .A(n62625), .ZN(n27208) );
  INV_X1 U31679 ( .A(n27208), .ZN(p_wishbone_bd_ram_n24408) );
  INV_X1 U31680 ( .A(n62624), .ZN(n27210) );
  INV_X1 U31681 ( .A(n27210), .ZN(p_wishbone_bd_ram_n24407) );
  INV_X1 U31682 ( .A(n62623), .ZN(n27212) );
  INV_X1 U31683 ( .A(n27212), .ZN(p_wishbone_bd_ram_n24406) );
  INV_X1 U31684 ( .A(n62622), .ZN(n27214) );
  INV_X1 U31685 ( .A(n27214), .ZN(p_wishbone_bd_ram_n24405) );
  INV_X1 U31686 ( .A(n62621), .ZN(n27216) );
  INV_X1 U31687 ( .A(n27216), .ZN(p_wishbone_bd_ram_n24404) );
  INV_X1 U31688 ( .A(n62620), .ZN(n27218) );
  INV_X1 U31689 ( .A(n27218), .ZN(p_wishbone_bd_ram_n24403) );
  INV_X1 U31690 ( .A(n62619), .ZN(n27220) );
  INV_X1 U31691 ( .A(n27220), .ZN(p_wishbone_bd_ram_n24402) );
  INV_X1 U31692 ( .A(n62618), .ZN(n27222) );
  INV_X1 U31693 ( .A(n27222), .ZN(p_wishbone_bd_ram_n24401) );
  INV_X1 U31694 ( .A(n62617), .ZN(n27224) );
  INV_X1 U31695 ( .A(n27224), .ZN(p_wishbone_bd_ram_n24400) );
  INV_X1 U31696 ( .A(n62616), .ZN(n27226) );
  INV_X1 U31697 ( .A(n27226), .ZN(p_wishbone_bd_ram_n24399) );
  INV_X1 U31698 ( .A(n62615), .ZN(n27228) );
  INV_X1 U31699 ( .A(n27228), .ZN(p_wishbone_bd_ram_n24398) );
  INV_X1 U31700 ( .A(n62614), .ZN(n27230) );
  INV_X1 U31701 ( .A(n27230), .ZN(p_wishbone_bd_ram_n24397) );
  INV_X1 U31702 ( .A(n62613), .ZN(n27232) );
  INV_X1 U31703 ( .A(n27232), .ZN(p_wishbone_bd_ram_n24396) );
  INV_X1 U31704 ( .A(n62612), .ZN(n27234) );
  INV_X1 U31705 ( .A(n27234), .ZN(p_wishbone_bd_ram_n24395) );
  INV_X1 U31706 ( .A(n62611), .ZN(n27236) );
  INV_X1 U31707 ( .A(n27236), .ZN(p_wishbone_bd_ram_n24394) );
  INV_X1 U31708 ( .A(n62610), .ZN(n27238) );
  INV_X1 U31709 ( .A(n27238), .ZN(p_wishbone_bd_ram_n24393) );
  INV_X1 U31710 ( .A(n62609), .ZN(n27240) );
  INV_X1 U31711 ( .A(n27240), .ZN(p_wishbone_bd_ram_n24392) );
  INV_X1 U31712 ( .A(n62608), .ZN(n27242) );
  INV_X1 U31713 ( .A(n27242), .ZN(p_wishbone_bd_ram_n24391) );
  INV_X1 U31714 ( .A(n62607), .ZN(n27244) );
  INV_X1 U31715 ( .A(n27244), .ZN(p_wishbone_bd_ram_n24390) );
  INV_X1 U31716 ( .A(n62606), .ZN(n27246) );
  INV_X1 U31717 ( .A(n27246), .ZN(p_wishbone_bd_ram_n24389) );
  INV_X1 U31718 ( .A(n62605), .ZN(n27248) );
  INV_X1 U31719 ( .A(n27248), .ZN(p_wishbone_bd_ram_n24388) );
  INV_X1 U31720 ( .A(n62604), .ZN(n27250) );
  INV_X1 U31721 ( .A(n27250), .ZN(p_wishbone_bd_ram_n24387) );
  INV_X1 U31722 ( .A(n62603), .ZN(n27252) );
  INV_X1 U31723 ( .A(n27252), .ZN(p_wishbone_bd_ram_n24386) );
  INV_X1 U31724 ( .A(n62602), .ZN(n27254) );
  INV_X1 U31725 ( .A(n27254), .ZN(p_wishbone_bd_ram_n24385) );
  INV_X1 U31726 ( .A(n62601), .ZN(n27256) );
  INV_X1 U31727 ( .A(n27256), .ZN(p_wishbone_bd_ram_n24384) );
  INV_X1 U31728 ( .A(n62600), .ZN(n27258) );
  INV_X1 U31729 ( .A(n27258), .ZN(p_wishbone_bd_ram_n24383) );
  INV_X1 U31730 ( .A(n62599), .ZN(n27260) );
  INV_X1 U31731 ( .A(n27260), .ZN(p_wishbone_bd_ram_n24382) );
  INV_X1 U31732 ( .A(n62598), .ZN(n27262) );
  INV_X1 U31733 ( .A(n27262), .ZN(p_wishbone_bd_ram_n24381) );
  INV_X1 U31734 ( .A(n62597), .ZN(n27264) );
  INV_X1 U31735 ( .A(n27264), .ZN(p_wishbone_bd_ram_n24380) );
  INV_X1 U31736 ( .A(n62596), .ZN(n27266) );
  INV_X1 U31737 ( .A(n27266), .ZN(p_wishbone_bd_ram_n24379) );
  INV_X1 U31738 ( .A(n62595), .ZN(n27268) );
  INV_X1 U31739 ( .A(n27268), .ZN(p_wishbone_bd_ram_n24378) );
  INV_X1 U31740 ( .A(n62594), .ZN(n27270) );
  INV_X1 U31741 ( .A(n27270), .ZN(p_wishbone_bd_ram_n24377) );
  INV_X1 U31742 ( .A(n62593), .ZN(n27272) );
  INV_X1 U31743 ( .A(n27272), .ZN(p_wishbone_bd_ram_n24376) );
  INV_X1 U31744 ( .A(n62592), .ZN(n27274) );
  INV_X1 U31745 ( .A(n27274), .ZN(p_wishbone_bd_ram_n24375) );
  INV_X1 U31746 ( .A(n62591), .ZN(n27276) );
  INV_X1 U31747 ( .A(n27276), .ZN(p_wishbone_bd_ram_n24374) );
  INV_X1 U31748 ( .A(n62590), .ZN(n27278) );
  INV_X1 U31749 ( .A(n27278), .ZN(p_wishbone_bd_ram_n24373) );
  INV_X1 U31750 ( .A(n62589), .ZN(n27280) );
  INV_X1 U31751 ( .A(n27280), .ZN(p_wishbone_bd_ram_n24372) );
  INV_X1 U31752 ( .A(n62588), .ZN(n27282) );
  INV_X1 U31753 ( .A(n27282), .ZN(p_wishbone_bd_ram_n24371) );
  INV_X1 U31754 ( .A(n62587), .ZN(n27284) );
  INV_X1 U31755 ( .A(n27284), .ZN(p_wishbone_bd_ram_n24370) );
  INV_X1 U31756 ( .A(n62586), .ZN(n27286) );
  INV_X1 U31757 ( .A(n27286), .ZN(p_wishbone_bd_ram_n24369) );
  INV_X1 U31758 ( .A(n62585), .ZN(n27288) );
  INV_X1 U31759 ( .A(n27288), .ZN(p_wishbone_bd_ram_n24367) );
  INV_X1 U31760 ( .A(n62584), .ZN(n27290) );
  INV_X1 U31761 ( .A(n27290), .ZN(p_wishbone_bd_ram_n24365) );
  INV_X1 U31762 ( .A(n62583), .ZN(n27292) );
  INV_X1 U31763 ( .A(n27292), .ZN(p_wishbone_bd_ram_n24364) );
  INV_X1 U31764 ( .A(n62582), .ZN(n27294) );
  INV_X1 U31765 ( .A(n27294), .ZN(p_wishbone_bd_ram_n24362) );
  INV_X1 U31766 ( .A(n62581), .ZN(n27296) );
  INV_X1 U31767 ( .A(n27296), .ZN(p_wishbone_bd_ram_n24360) );
  INV_X1 U31768 ( .A(n62580), .ZN(n27298) );
  INV_X1 U31769 ( .A(n27298), .ZN(p_wishbone_bd_ram_n24359) );
  INV_X1 U31770 ( .A(n62579), .ZN(n27300) );
  INV_X1 U31771 ( .A(n27300), .ZN(p_wishbone_bd_ram_n24358) );
  INV_X1 U31772 ( .A(n62578), .ZN(n27302) );
  INV_X1 U31773 ( .A(n27302), .ZN(p_wishbone_bd_ram_n24357) );
  INV_X1 U31774 ( .A(n62577), .ZN(n27304) );
  INV_X1 U31775 ( .A(n27304), .ZN(p_wishbone_bd_ram_n24356) );
  INV_X1 U31776 ( .A(n62576), .ZN(n27306) );
  INV_X1 U31777 ( .A(n27306), .ZN(p_wishbone_bd_ram_n24355) );
  INV_X1 U31778 ( .A(n62575), .ZN(n27308) );
  INV_X1 U31779 ( .A(n27308), .ZN(p_wishbone_bd_ram_n24354) );
  INV_X1 U31780 ( .A(n62574), .ZN(n27310) );
  INV_X1 U31781 ( .A(n27310), .ZN(p_wishbone_bd_ram_n24353) );
  INV_X1 U31782 ( .A(n62573), .ZN(n27312) );
  INV_X1 U31783 ( .A(n27312), .ZN(p_wishbone_bd_ram_n24352) );
  INV_X1 U31784 ( .A(n62572), .ZN(n27314) );
  INV_X1 U31785 ( .A(n27314), .ZN(p_wishbone_bd_ram_n24350) );
  INV_X1 U31786 ( .A(n62571), .ZN(n27316) );
  INV_X1 U31787 ( .A(n27316), .ZN(p_wishbone_bd_ram_n24347) );
  INV_X1 U31788 ( .A(n62570), .ZN(n27318) );
  INV_X1 U31789 ( .A(n27318), .ZN(p_wishbone_bd_ram_n24345) );
  INV_X1 U31790 ( .A(n62569), .ZN(n27320) );
  INV_X1 U31791 ( .A(n27320), .ZN(p_wishbone_bd_ram_n24344) );
  INV_X1 U31792 ( .A(n62568), .ZN(n27322) );
  INV_X1 U31793 ( .A(n27322), .ZN(p_wishbone_bd_ram_n24343) );
  INV_X1 U31794 ( .A(n62567), .ZN(n27324) );
  INV_X1 U31795 ( .A(n27324), .ZN(p_wishbone_bd_ram_n24342) );
  INV_X1 U31796 ( .A(n62566), .ZN(n27326) );
  INV_X1 U31797 ( .A(n27326), .ZN(p_wishbone_bd_ram_n24341) );
  INV_X1 U31798 ( .A(n62565), .ZN(n27328) );
  INV_X1 U31799 ( .A(n27328), .ZN(p_wishbone_bd_ram_n24340) );
  INV_X1 U31800 ( .A(n62564), .ZN(n27330) );
  INV_X1 U31801 ( .A(n27330), .ZN(p_wishbone_bd_ram_n24339) );
  INV_X1 U31802 ( .A(n62563), .ZN(n27332) );
  INV_X1 U31803 ( .A(n27332), .ZN(p_wishbone_bd_ram_n24338) );
  INV_X1 U31804 ( .A(n62562), .ZN(n27334) );
  INV_X1 U31805 ( .A(n27334), .ZN(p_wishbone_bd_ram_n24337) );
  INV_X1 U31806 ( .A(n62561), .ZN(n27336) );
  INV_X1 U31807 ( .A(n27336), .ZN(p_wishbone_bd_ram_n24336) );
  INV_X1 U31808 ( .A(n62560), .ZN(n27338) );
  INV_X1 U31809 ( .A(n27338), .ZN(p_wishbone_bd_ram_n24335) );
  INV_X1 U31810 ( .A(n62559), .ZN(n27340) );
  INV_X1 U31811 ( .A(n27340), .ZN(p_wishbone_bd_ram_n24334) );
  INV_X1 U31812 ( .A(n62558), .ZN(n27342) );
  INV_X1 U31813 ( .A(n27342), .ZN(p_wishbone_bd_ram_n24333) );
  INV_X1 U31814 ( .A(n62557), .ZN(n27344) );
  INV_X1 U31815 ( .A(n27344), .ZN(p_wishbone_bd_ram_n24332) );
  INV_X1 U31816 ( .A(n62556), .ZN(n27346) );
  INV_X1 U31817 ( .A(n27346), .ZN(p_wishbone_bd_ram_n24331) );
  INV_X1 U31818 ( .A(n62555), .ZN(n27348) );
  INV_X1 U31819 ( .A(n27348), .ZN(p_wishbone_bd_ram_n24330) );
  INV_X1 U31820 ( .A(n62554), .ZN(n27350) );
  INV_X1 U31821 ( .A(n27350), .ZN(p_wishbone_bd_ram_n24329) );
  INV_X1 U31822 ( .A(n62553), .ZN(n27352) );
  INV_X1 U31823 ( .A(n27352), .ZN(p_wishbone_bd_ram_n24328) );
  INV_X1 U31824 ( .A(n62552), .ZN(n27354) );
  INV_X1 U31825 ( .A(n27354), .ZN(p_wishbone_bd_ram_n24327) );
  INV_X1 U31826 ( .A(n62551), .ZN(n27356) );
  INV_X1 U31827 ( .A(n27356), .ZN(p_wishbone_bd_ram_n24326) );
  INV_X1 U31828 ( .A(n62550), .ZN(n27358) );
  INV_X1 U31829 ( .A(n27358), .ZN(p_wishbone_bd_ram_n24325) );
  INV_X1 U31830 ( .A(n62549), .ZN(n27360) );
  INV_X1 U31831 ( .A(n27360), .ZN(p_wishbone_bd_ram_n24324) );
  INV_X1 U31832 ( .A(n62548), .ZN(n27362) );
  INV_X1 U31833 ( .A(n27362), .ZN(p_wishbone_bd_ram_n24323) );
  INV_X1 U31834 ( .A(n62547), .ZN(n27364) );
  INV_X1 U31835 ( .A(n27364), .ZN(p_wishbone_bd_ram_n24322) );
  INV_X1 U31836 ( .A(n62546), .ZN(n27366) );
  INV_X1 U31837 ( .A(n27366), .ZN(p_wishbone_bd_ram_n24321) );
  INV_X1 U31838 ( .A(n62545), .ZN(n27368) );
  INV_X1 U31839 ( .A(n27368), .ZN(p_wishbone_bd_ram_n24320) );
  INV_X1 U31840 ( .A(n62544), .ZN(n27370) );
  INV_X1 U31841 ( .A(n27370), .ZN(p_wishbone_bd_ram_n24319) );
  INV_X1 U31842 ( .A(n62543), .ZN(n27372) );
  INV_X1 U31843 ( .A(n27372), .ZN(p_wishbone_bd_ram_n24318) );
  INV_X1 U31844 ( .A(n62542), .ZN(n27374) );
  INV_X1 U31845 ( .A(n27374), .ZN(p_wishbone_bd_ram_n24317) );
  INV_X1 U31846 ( .A(n62541), .ZN(n27376) );
  INV_X1 U31847 ( .A(n27376), .ZN(p_wishbone_bd_ram_n24316) );
  INV_X1 U31848 ( .A(n62540), .ZN(n27378) );
  INV_X1 U31849 ( .A(n27378), .ZN(p_wishbone_bd_ram_n24315) );
  INV_X1 U31850 ( .A(n62539), .ZN(n27380) );
  INV_X1 U31851 ( .A(n27380), .ZN(p_wishbone_bd_ram_n24314) );
  INV_X1 U31852 ( .A(n62538), .ZN(n27382) );
  INV_X1 U31853 ( .A(n27382), .ZN(p_wishbone_bd_ram_n24313) );
  INV_X1 U31854 ( .A(n62537), .ZN(n27384) );
  INV_X1 U31855 ( .A(n27384), .ZN(p_wishbone_bd_ram_n24312) );
  INV_X1 U31856 ( .A(n62536), .ZN(n27386) );
  INV_X1 U31857 ( .A(n27386), .ZN(p_wishbone_bd_ram_n24311) );
  INV_X1 U31858 ( .A(n62535), .ZN(n27388) );
  INV_X1 U31859 ( .A(n27388), .ZN(p_wishbone_bd_ram_n24310) );
  INV_X1 U31860 ( .A(n62534), .ZN(n27390) );
  INV_X1 U31861 ( .A(n27390), .ZN(p_wishbone_bd_ram_n24309) );
  INV_X1 U31862 ( .A(n62533), .ZN(n27392) );
  INV_X1 U31863 ( .A(n27392), .ZN(p_wishbone_bd_ram_n24308) );
  INV_X1 U31864 ( .A(n62532), .ZN(n27394) );
  INV_X1 U31865 ( .A(n27394), .ZN(p_wishbone_bd_ram_n24307) );
  INV_X1 U31866 ( .A(n62531), .ZN(n27396) );
  INV_X1 U31867 ( .A(n27396), .ZN(p_wishbone_bd_ram_n24306) );
  INV_X1 U31868 ( .A(n62530), .ZN(n27398) );
  INV_X1 U31869 ( .A(n27398), .ZN(p_wishbone_bd_ram_n24305) );
  INV_X1 U31870 ( .A(n62529), .ZN(n27400) );
  INV_X1 U31871 ( .A(n27400), .ZN(p_wishbone_bd_ram_n24304) );
  INV_X1 U31872 ( .A(n62528), .ZN(n27402) );
  INV_X1 U31873 ( .A(n27402), .ZN(p_wishbone_bd_ram_n24303) );
  INV_X1 U31874 ( .A(n62527), .ZN(n27404) );
  INV_X1 U31875 ( .A(n27404), .ZN(p_wishbone_bd_ram_n24302) );
  INV_X1 U31876 ( .A(n62526), .ZN(n27406) );
  INV_X1 U31877 ( .A(n27406), .ZN(p_wishbone_bd_ram_n24301) );
  INV_X1 U31878 ( .A(n62525), .ZN(n27408) );
  INV_X1 U31879 ( .A(n27408), .ZN(p_wishbone_bd_ram_n24300) );
  INV_X1 U31880 ( .A(n62524), .ZN(n27410) );
  INV_X1 U31881 ( .A(n27410), .ZN(p_wishbone_bd_ram_n24299) );
  INV_X1 U31882 ( .A(n62523), .ZN(n27412) );
  INV_X1 U31883 ( .A(n27412), .ZN(p_wishbone_bd_ram_n24298) );
  INV_X1 U31884 ( .A(n62522), .ZN(n27414) );
  INV_X1 U31885 ( .A(n27414), .ZN(p_wishbone_bd_ram_n24297) );
  INV_X1 U31886 ( .A(n62521), .ZN(n27416) );
  INV_X1 U31887 ( .A(n27416), .ZN(p_wishbone_bd_ram_n24296) );
  INV_X1 U31888 ( .A(n62520), .ZN(n27418) );
  INV_X1 U31889 ( .A(n27418), .ZN(p_wishbone_bd_ram_n24294) );
  INV_X1 U31890 ( .A(n62519), .ZN(n27420) );
  INV_X1 U31891 ( .A(n27420), .ZN(p_wishbone_bd_ram_n24291) );
  INV_X1 U31892 ( .A(n62518), .ZN(n27422) );
  INV_X1 U31893 ( .A(n27422), .ZN(p_wishbone_bd_ram_n24289) );
  INV_X1 U31894 ( .A(n62517), .ZN(n27424) );
  INV_X1 U31895 ( .A(n27424), .ZN(p_wishbone_bd_ram_n24288) );
  INV_X1 U31896 ( .A(n62516), .ZN(n27426) );
  INV_X1 U31897 ( .A(n27426), .ZN(p_wishbone_bd_ram_n24287) );
  INV_X1 U31898 ( .A(n62515), .ZN(n27428) );
  INV_X1 U31899 ( .A(n27428), .ZN(p_wishbone_bd_ram_n24286) );
  INV_X1 U31900 ( .A(n62514), .ZN(n27430) );
  INV_X1 U31901 ( .A(n27430), .ZN(p_wishbone_bd_ram_n24285) );
  INV_X1 U31902 ( .A(n62513), .ZN(n27432) );
  INV_X1 U31903 ( .A(n27432), .ZN(p_wishbone_bd_ram_n24284) );
  INV_X1 U31904 ( .A(n62512), .ZN(n27434) );
  INV_X1 U31905 ( .A(n27434), .ZN(p_wishbone_bd_ram_n24283) );
  INV_X1 U31906 ( .A(n62511), .ZN(n27436) );
  INV_X1 U31907 ( .A(n27436), .ZN(p_wishbone_bd_ram_n24282) );
  INV_X1 U31908 ( .A(n62510), .ZN(n27438) );
  INV_X1 U31909 ( .A(n27438), .ZN(p_wishbone_bd_ram_n24281) );
  INV_X1 U31910 ( .A(n62509), .ZN(n27440) );
  INV_X1 U31911 ( .A(n27440), .ZN(p_wishbone_bd_ram_n24280) );
  INV_X1 U31912 ( .A(n62508), .ZN(n27442) );
  INV_X1 U31913 ( .A(n27442), .ZN(p_wishbone_bd_ram_n24279) );
  INV_X1 U31914 ( .A(n62507), .ZN(n27444) );
  INV_X1 U31915 ( .A(n27444), .ZN(p_wishbone_bd_ram_n24278) );
  INV_X1 U31916 ( .A(n62506), .ZN(n27446) );
  INV_X1 U31917 ( .A(n27446), .ZN(p_wishbone_bd_ram_n24277) );
  INV_X1 U31918 ( .A(n62505), .ZN(n27448) );
  INV_X1 U31919 ( .A(n27448), .ZN(p_wishbone_bd_ram_n24276) );
  INV_X1 U31920 ( .A(n62504), .ZN(n27450) );
  INV_X1 U31921 ( .A(n27450), .ZN(p_wishbone_bd_ram_n24275) );
  INV_X1 U31922 ( .A(n62503), .ZN(n27452) );
  INV_X1 U31923 ( .A(n27452), .ZN(p_wishbone_bd_ram_n24274) );
  INV_X1 U31924 ( .A(n62502), .ZN(n27454) );
  INV_X1 U31925 ( .A(n27454), .ZN(p_wishbone_bd_ram_n24273) );
  INV_X1 U31926 ( .A(n62501), .ZN(n27456) );
  INV_X1 U31927 ( .A(n27456), .ZN(p_wishbone_bd_ram_n24272) );
  INV_X1 U31928 ( .A(n62500), .ZN(n27458) );
  INV_X1 U31929 ( .A(n27458), .ZN(p_wishbone_bd_ram_n24271) );
  INV_X1 U31930 ( .A(n62499), .ZN(n27460) );
  INV_X1 U31931 ( .A(n27460), .ZN(p_wishbone_bd_ram_n24270) );
  INV_X1 U31932 ( .A(n62498), .ZN(n27462) );
  INV_X1 U31933 ( .A(n27462), .ZN(p_wishbone_bd_ram_n24269) );
  INV_X1 U31934 ( .A(n62497), .ZN(n27464) );
  INV_X1 U31935 ( .A(n27464), .ZN(p_wishbone_bd_ram_n24268) );
  INV_X1 U31936 ( .A(n62496), .ZN(n27466) );
  INV_X1 U31937 ( .A(n27466), .ZN(p_wishbone_bd_ram_n24267) );
  INV_X1 U31938 ( .A(n62495), .ZN(n27468) );
  INV_X1 U31939 ( .A(n27468), .ZN(p_wishbone_bd_ram_n24266) );
  INV_X1 U31940 ( .A(n62494), .ZN(n27470) );
  INV_X1 U31941 ( .A(n27470), .ZN(p_wishbone_bd_ram_n24265) );
  INV_X1 U31942 ( .A(n62493), .ZN(n27472) );
  INV_X1 U31943 ( .A(n27472), .ZN(p_wishbone_bd_ram_n24263) );
  INV_X1 U31944 ( .A(n62492), .ZN(n27474) );
  INV_X1 U31945 ( .A(n27474), .ZN(p_wishbone_bd_ram_n24261) );
  INV_X1 U31946 ( .A(n62491), .ZN(n27476) );
  INV_X1 U31947 ( .A(n27476), .ZN(p_wishbone_bd_ram_n24260) );
  INV_X1 U31948 ( .A(n62490), .ZN(n27478) );
  INV_X1 U31949 ( .A(n27478), .ZN(p_wishbone_bd_ram_n24258) );
  INV_X1 U31950 ( .A(n62489), .ZN(n27480) );
  INV_X1 U31951 ( .A(n27480), .ZN(p_wishbone_bd_ram_n24256) );
  INV_X1 U31952 ( .A(n62488), .ZN(n27482) );
  INV_X1 U31953 ( .A(n27482), .ZN(p_wishbone_bd_ram_n24255) );
  INV_X1 U31954 ( .A(n62487), .ZN(n27484) );
  INV_X1 U31955 ( .A(n27484), .ZN(p_wishbone_bd_ram_n24254) );
  INV_X1 U31956 ( .A(n62486), .ZN(n27486) );
  INV_X1 U31957 ( .A(n27486), .ZN(p_wishbone_bd_ram_n24253) );
  INV_X1 U31958 ( .A(n62485), .ZN(n27488) );
  INV_X1 U31959 ( .A(n27488), .ZN(p_wishbone_bd_ram_n24252) );
  INV_X1 U31960 ( .A(n62484), .ZN(n27490) );
  INV_X1 U31961 ( .A(n27490), .ZN(p_wishbone_bd_ram_n24251) );
  INV_X1 U31962 ( .A(n62483), .ZN(n27492) );
  INV_X1 U31963 ( .A(n27492), .ZN(p_wishbone_bd_ram_n24250) );
  INV_X1 U31964 ( .A(n62482), .ZN(n27494) );
  INV_X1 U31965 ( .A(n27494), .ZN(p_wishbone_bd_ram_n24249) );
  INV_X1 U31966 ( .A(n62481), .ZN(n27496) );
  INV_X1 U31967 ( .A(n27496), .ZN(p_wishbone_bd_ram_n24248) );
  INV_X1 U31968 ( .A(n62480), .ZN(n27498) );
  INV_X1 U31969 ( .A(n27498), .ZN(p_wishbone_bd_ram_n24247) );
  INV_X1 U31970 ( .A(n62479), .ZN(n27500) );
  INV_X1 U31971 ( .A(n27500), .ZN(p_wishbone_bd_ram_n24246) );
  INV_X1 U31972 ( .A(n62478), .ZN(n27502) );
  INV_X1 U31973 ( .A(n27502), .ZN(p_wishbone_bd_ram_n24245) );
  INV_X1 U31974 ( .A(n62477), .ZN(n27504) );
  INV_X1 U31975 ( .A(n27504), .ZN(p_wishbone_bd_ram_n24244) );
  INV_X1 U31976 ( .A(n62476), .ZN(n27506) );
  INV_X1 U31977 ( .A(n27506), .ZN(p_wishbone_bd_ram_n24243) );
  INV_X1 U31978 ( .A(n62475), .ZN(n27508) );
  INV_X1 U31979 ( .A(n27508), .ZN(p_wishbone_bd_ram_n24242) );
  INV_X1 U31980 ( .A(n62474), .ZN(n27510) );
  INV_X1 U31981 ( .A(n27510), .ZN(p_wishbone_bd_ram_n24241) );
  INV_X1 U31982 ( .A(n62473), .ZN(n27512) );
  INV_X1 U31983 ( .A(n27512), .ZN(p_wishbone_bd_ram_n24240) );
  INV_X1 U31984 ( .A(n62472), .ZN(n27514) );
  INV_X1 U31985 ( .A(n27514), .ZN(p_wishbone_bd_ram_n24239) );
  INV_X1 U31986 ( .A(n62471), .ZN(n27516) );
  INV_X1 U31987 ( .A(n27516), .ZN(p_wishbone_bd_ram_n24238) );
  INV_X1 U31988 ( .A(n62470), .ZN(n27518) );
  INV_X1 U31989 ( .A(n27518), .ZN(p_wishbone_bd_ram_n24237) );
  INV_X1 U31990 ( .A(n62469), .ZN(n27520) );
  INV_X1 U31991 ( .A(n27520), .ZN(p_wishbone_bd_ram_n24236) );
  INV_X1 U31992 ( .A(n62468), .ZN(n27522) );
  INV_X1 U31993 ( .A(n27522), .ZN(p_wishbone_bd_ram_n24235) );
  INV_X1 U31994 ( .A(n62467), .ZN(n27524) );
  INV_X1 U31995 ( .A(n27524), .ZN(p_wishbone_bd_ram_n24234) );
  INV_X1 U31996 ( .A(n62466), .ZN(n27526) );
  INV_X1 U31997 ( .A(n27526), .ZN(p_wishbone_bd_ram_n24233) );
  INV_X1 U31998 ( .A(n62465), .ZN(n27528) );
  INV_X1 U31999 ( .A(n27528), .ZN(p_wishbone_bd_ram_n24232) );
  INV_X1 U32000 ( .A(n62464), .ZN(n27530) );
  INV_X1 U32001 ( .A(n27530), .ZN(p_wishbone_bd_ram_n24231) );
  INV_X1 U32002 ( .A(n62463), .ZN(n27532) );
  INV_X1 U32003 ( .A(n27532), .ZN(p_wishbone_bd_ram_n24230) );
  INV_X1 U32004 ( .A(n62462), .ZN(n27534) );
  INV_X1 U32005 ( .A(n27534), .ZN(p_wishbone_bd_ram_n24229) );
  INV_X1 U32006 ( .A(n62461), .ZN(n27536) );
  INV_X1 U32007 ( .A(n27536), .ZN(p_wishbone_bd_ram_n24228) );
  INV_X1 U32008 ( .A(n62460), .ZN(n27538) );
  INV_X1 U32009 ( .A(n27538), .ZN(p_wishbone_bd_ram_n24227) );
  INV_X1 U32010 ( .A(n62459), .ZN(n27540) );
  INV_X1 U32011 ( .A(n27540), .ZN(p_wishbone_bd_ram_n24226) );
  INV_X1 U32012 ( .A(n62458), .ZN(n27542) );
  INV_X1 U32013 ( .A(n27542), .ZN(p_wishbone_bd_ram_n24225) );
  INV_X1 U32014 ( .A(n62457), .ZN(n27544) );
  INV_X1 U32015 ( .A(n27544), .ZN(p_wishbone_bd_ram_n24224) );
  INV_X1 U32016 ( .A(n62456), .ZN(n27546) );
  INV_X1 U32017 ( .A(n27546), .ZN(p_wishbone_bd_ram_n24223) );
  INV_X1 U32018 ( .A(n62455), .ZN(n27548) );
  INV_X1 U32019 ( .A(n27548), .ZN(p_wishbone_bd_ram_n24222) );
  INV_X1 U32020 ( .A(n62454), .ZN(n27550) );
  INV_X1 U32021 ( .A(n27550), .ZN(p_wishbone_bd_ram_n24221) );
  INV_X1 U32022 ( .A(n62453), .ZN(n27552) );
  INV_X1 U32023 ( .A(n27552), .ZN(p_wishbone_bd_ram_n24220) );
  INV_X1 U32024 ( .A(n62452), .ZN(n27554) );
  INV_X1 U32025 ( .A(n27554), .ZN(p_wishbone_bd_ram_n24219) );
  INV_X1 U32026 ( .A(n62451), .ZN(n27556) );
  INV_X1 U32027 ( .A(n27556), .ZN(p_wishbone_bd_ram_n24218) );
  INV_X1 U32028 ( .A(n62450), .ZN(n27558) );
  INV_X1 U32029 ( .A(n27558), .ZN(p_wishbone_bd_ram_n24217) );
  INV_X1 U32030 ( .A(n62449), .ZN(n27560) );
  INV_X1 U32031 ( .A(n27560), .ZN(p_wishbone_bd_ram_n24216) );
  INV_X1 U32032 ( .A(n62448), .ZN(n27562) );
  INV_X1 U32033 ( .A(n27562), .ZN(p_wishbone_bd_ram_n24215) );
  INV_X1 U32034 ( .A(n62447), .ZN(n27564) );
  INV_X1 U32035 ( .A(n27564), .ZN(p_wishbone_bd_ram_n24214) );
  INV_X1 U32036 ( .A(n62446), .ZN(n27566) );
  INV_X1 U32037 ( .A(n27566), .ZN(p_wishbone_bd_ram_n24213) );
  INV_X1 U32038 ( .A(n62445), .ZN(n27568) );
  INV_X1 U32039 ( .A(n27568), .ZN(p_wishbone_bd_ram_n24212) );
  INV_X1 U32040 ( .A(n62444), .ZN(n27570) );
  INV_X1 U32041 ( .A(n27570), .ZN(p_wishbone_bd_ram_n24211) );
  INV_X1 U32042 ( .A(n62443), .ZN(n27572) );
  INV_X1 U32043 ( .A(n27572), .ZN(p_wishbone_bd_ram_n24210) );
  INV_X1 U32044 ( .A(n62442), .ZN(n27574) );
  INV_X1 U32045 ( .A(n27574), .ZN(p_wishbone_bd_ram_n24209) );
  INV_X1 U32046 ( .A(n62441), .ZN(n27576) );
  INV_X1 U32047 ( .A(n27576), .ZN(p_wishbone_bd_ram_n24208) );
  INV_X1 U32048 ( .A(n62440), .ZN(n27578) );
  INV_X1 U32049 ( .A(n27578), .ZN(p_wishbone_bd_ram_n24207) );
  INV_X1 U32050 ( .A(n62439), .ZN(n27580) );
  INV_X1 U32051 ( .A(n27580), .ZN(p_wishbone_bd_ram_n24206) );
  INV_X1 U32052 ( .A(n62438), .ZN(n27582) );
  INV_X1 U32053 ( .A(n27582), .ZN(p_wishbone_bd_ram_n24205) );
  INV_X1 U32054 ( .A(n62437), .ZN(n27584) );
  INV_X1 U32055 ( .A(n27584), .ZN(p_wishbone_bd_ram_n24204) );
  INV_X1 U32056 ( .A(n62436), .ZN(n27586) );
  INV_X1 U32057 ( .A(n27586), .ZN(p_wishbone_bd_ram_n24203) );
  INV_X1 U32058 ( .A(n62435), .ZN(n27588) );
  INV_X1 U32059 ( .A(n27588), .ZN(p_wishbone_bd_ram_n24202) );
  INV_X1 U32060 ( .A(n62434), .ZN(n27590) );
  INV_X1 U32061 ( .A(n27590), .ZN(p_wishbone_bd_ram_n24201) );
  INV_X1 U32062 ( .A(n62433), .ZN(n27592) );
  INV_X1 U32063 ( .A(n27592), .ZN(p_wishbone_bd_ram_n24200) );
  INV_X1 U32064 ( .A(n62432), .ZN(n27594) );
  INV_X1 U32065 ( .A(n27594), .ZN(p_wishbone_bd_ram_n24198) );
  INV_X1 U32066 ( .A(n62431), .ZN(n27596) );
  INV_X1 U32067 ( .A(n27596), .ZN(p_wishbone_bd_ram_n24195) );
  INV_X1 U32068 ( .A(n62430), .ZN(n27598) );
  INV_X1 U32069 ( .A(n27598), .ZN(p_wishbone_bd_ram_n24193) );
  INV_X1 U32070 ( .A(n62429), .ZN(n27600) );
  INV_X1 U32071 ( .A(n27600), .ZN(p_wishbone_bd_ram_n24192) );
  INV_X1 U32072 ( .A(n62428), .ZN(n27602) );
  INV_X1 U32073 ( .A(n27602), .ZN(p_wishbone_bd_ram_n24191) );
  INV_X1 U32074 ( .A(n62427), .ZN(n27604) );
  INV_X1 U32075 ( .A(n27604), .ZN(p_wishbone_bd_ram_n24190) );
  INV_X1 U32076 ( .A(n62426), .ZN(n27606) );
  INV_X1 U32077 ( .A(n27606), .ZN(p_wishbone_bd_ram_n24189) );
  INV_X1 U32078 ( .A(n62425), .ZN(n27608) );
  INV_X1 U32079 ( .A(n27608), .ZN(p_wishbone_bd_ram_n24188) );
  INV_X1 U32080 ( .A(n62424), .ZN(n27610) );
  INV_X1 U32081 ( .A(n27610), .ZN(p_wishbone_bd_ram_n24187) );
  INV_X1 U32082 ( .A(n62423), .ZN(n27612) );
  INV_X1 U32083 ( .A(n27612), .ZN(p_wishbone_bd_ram_n24186) );
  INV_X1 U32084 ( .A(n62422), .ZN(n27614) );
  INV_X1 U32085 ( .A(n27614), .ZN(p_wishbone_bd_ram_n24185) );
  INV_X1 U32086 ( .A(n62421), .ZN(n27616) );
  INV_X1 U32087 ( .A(n27616), .ZN(p_wishbone_bd_ram_n24183) );
  INV_X1 U32088 ( .A(n62420), .ZN(n27618) );
  INV_X1 U32089 ( .A(n27618), .ZN(p_wishbone_bd_ram_n24181) );
  INV_X1 U32090 ( .A(n62419), .ZN(n27620) );
  INV_X1 U32091 ( .A(n27620), .ZN(p_wishbone_bd_ram_n24180) );
  INV_X1 U32092 ( .A(n62418), .ZN(n27622) );
  INV_X1 U32093 ( .A(n27622), .ZN(p_wishbone_bd_ram_n24178) );
  INV_X1 U32094 ( .A(n62417), .ZN(n27624) );
  INV_X1 U32095 ( .A(n27624), .ZN(p_wishbone_bd_ram_n24175) );
  INV_X1 U32096 ( .A(n62416), .ZN(n27626) );
  INV_X1 U32097 ( .A(n27626), .ZN(p_wishbone_bd_ram_n24173) );
  INV_X1 U32098 ( .A(n62415), .ZN(n27628) );
  INV_X1 U32099 ( .A(n27628), .ZN(p_wishbone_bd_ram_n24172) );
  INV_X1 U32100 ( .A(n62414), .ZN(n27630) );
  INV_X1 U32101 ( .A(n27630), .ZN(p_wishbone_bd_ram_n24170) );
  INV_X1 U32102 ( .A(n62413), .ZN(n27632) );
  INV_X1 U32103 ( .A(n27632), .ZN(p_wishbone_bd_ram_n24167) );
  INV_X1 U32104 ( .A(n62412), .ZN(n27634) );
  INV_X1 U32105 ( .A(n27634), .ZN(p_wishbone_bd_ram_n24165) );
  INV_X1 U32106 ( .A(n62411), .ZN(n27636) );
  INV_X1 U32107 ( .A(n27636), .ZN(p_wishbone_bd_ram_n24164) );
  INV_X1 U32108 ( .A(n62410), .ZN(n27638) );
  INV_X1 U32109 ( .A(n27638), .ZN(p_wishbone_bd_ram_n24162) );
  INV_X1 U32110 ( .A(n62409), .ZN(n27640) );
  INV_X1 U32111 ( .A(n27640), .ZN(p_wishbone_bd_ram_n24160) );
  INV_X1 U32112 ( .A(n62408), .ZN(n27642) );
  INV_X1 U32113 ( .A(n27642), .ZN(p_wishbone_bd_ram_n24159) );
  INV_X1 U32114 ( .A(n62407), .ZN(n27644) );
  INV_X1 U32115 ( .A(n27644), .ZN(p_wishbone_bd_ram_n24158) );
  INV_X1 U32116 ( .A(n62406), .ZN(n27646) );
  INV_X1 U32117 ( .A(n27646), .ZN(p_wishbone_bd_ram_n24157) );
  INV_X1 U32118 ( .A(n62405), .ZN(n27648) );
  INV_X1 U32119 ( .A(n27648), .ZN(p_wishbone_bd_ram_n24156) );
  INV_X1 U32120 ( .A(n62404), .ZN(n27650) );
  INV_X1 U32121 ( .A(n27650), .ZN(p_wishbone_bd_ram_n24155) );
  INV_X1 U32122 ( .A(n62403), .ZN(n27652) );
  INV_X1 U32123 ( .A(n27652), .ZN(p_wishbone_bd_ram_n24154) );
  INV_X1 U32124 ( .A(n62402), .ZN(n27654) );
  INV_X1 U32125 ( .A(n27654), .ZN(p_wishbone_bd_ram_n24153) );
  INV_X1 U32126 ( .A(n62401), .ZN(n27656) );
  INV_X1 U32127 ( .A(n27656), .ZN(p_wishbone_bd_ram_n24152) );
  INV_X1 U32128 ( .A(n62400), .ZN(n27658) );
  INV_X1 U32129 ( .A(n27658), .ZN(p_wishbone_bd_ram_n24151) );
  INV_X1 U32130 ( .A(n62399), .ZN(n27660) );
  INV_X1 U32131 ( .A(n27660), .ZN(p_wishbone_bd_ram_n24150) );
  INV_X1 U32132 ( .A(n62398), .ZN(n27662) );
  INV_X1 U32133 ( .A(n27662), .ZN(p_wishbone_bd_ram_n24149) );
  INV_X1 U32134 ( .A(n62397), .ZN(n27664) );
  INV_X1 U32135 ( .A(n27664), .ZN(p_wishbone_bd_ram_n24148) );
  INV_X1 U32136 ( .A(n62396), .ZN(n27666) );
  INV_X1 U32137 ( .A(n27666), .ZN(p_wishbone_bd_ram_n24147) );
  INV_X1 U32138 ( .A(n62395), .ZN(n27668) );
  INV_X1 U32139 ( .A(n27668), .ZN(p_wishbone_bd_ram_n24146) );
  INV_X1 U32140 ( .A(n62394), .ZN(n27670) );
  INV_X1 U32141 ( .A(n27670), .ZN(p_wishbone_bd_ram_n24145) );
  INV_X1 U32142 ( .A(n62393), .ZN(n27672) );
  INV_X1 U32143 ( .A(n27672), .ZN(p_wishbone_bd_ram_n24144) );
  INV_X1 U32144 ( .A(n62392), .ZN(n27674) );
  INV_X1 U32145 ( .A(n27674), .ZN(p_wishbone_bd_ram_n24143) );
  INV_X1 U32146 ( .A(n62391), .ZN(n27676) );
  INV_X1 U32147 ( .A(n27676), .ZN(p_wishbone_bd_ram_n24142) );
  INV_X1 U32148 ( .A(n62390), .ZN(n27678) );
  INV_X1 U32149 ( .A(n27678), .ZN(p_wishbone_bd_ram_n24141) );
  INV_X1 U32150 ( .A(n62389), .ZN(n27680) );
  INV_X1 U32151 ( .A(n27680), .ZN(p_wishbone_bd_ram_n24140) );
  INV_X1 U32152 ( .A(n62388), .ZN(n27682) );
  INV_X1 U32153 ( .A(n27682), .ZN(p_wishbone_bd_ram_n24139) );
  INV_X1 U32154 ( .A(n62387), .ZN(n27684) );
  INV_X1 U32155 ( .A(n27684), .ZN(p_wishbone_bd_ram_n24138) );
  INV_X1 U32156 ( .A(n62386), .ZN(n27686) );
  INV_X1 U32157 ( .A(n27686), .ZN(p_wishbone_bd_ram_n24137) );
  INV_X1 U32158 ( .A(n62385), .ZN(n27688) );
  INV_X1 U32159 ( .A(n27688), .ZN(p_wishbone_bd_ram_n24135) );
  INV_X1 U32160 ( .A(n62384), .ZN(n27690) );
  INV_X1 U32161 ( .A(n27690), .ZN(p_wishbone_bd_ram_n24133) );
  INV_X1 U32162 ( .A(n62383), .ZN(n27692) );
  INV_X1 U32163 ( .A(n27692), .ZN(p_wishbone_bd_ram_n24132) );
  INV_X1 U32164 ( .A(n62382), .ZN(n27694) );
  INV_X1 U32165 ( .A(n27694), .ZN(p_wishbone_bd_ram_n24130) );
  INV_X1 U32166 ( .A(n62381), .ZN(n27696) );
  INV_X1 U32167 ( .A(n27696), .ZN(p_wishbone_bd_ram_n24128) );
  INV_X1 U32168 ( .A(n62380), .ZN(n27698) );
  INV_X1 U32169 ( .A(n27698), .ZN(p_wishbone_bd_ram_n24127) );
  INV_X1 U32170 ( .A(n62379), .ZN(n27700) );
  INV_X1 U32171 ( .A(n27700), .ZN(p_wishbone_bd_ram_n24126) );
  INV_X1 U32172 ( .A(n62378), .ZN(n27702) );
  INV_X1 U32173 ( .A(n27702), .ZN(p_wishbone_bd_ram_n24125) );
  INV_X1 U32174 ( .A(n62377), .ZN(n27704) );
  INV_X1 U32175 ( .A(n27704), .ZN(p_wishbone_bd_ram_n24124) );
  INV_X1 U32176 ( .A(n62376), .ZN(n27706) );
  INV_X1 U32177 ( .A(n27706), .ZN(p_wishbone_bd_ram_n24123) );
  INV_X1 U32178 ( .A(n62375), .ZN(n27708) );
  INV_X1 U32179 ( .A(n27708), .ZN(p_wishbone_bd_ram_n24122) );
  INV_X1 U32180 ( .A(n62374), .ZN(n27710) );
  INV_X1 U32181 ( .A(n27710), .ZN(p_wishbone_bd_ram_n24121) );
  INV_X1 U32182 ( .A(n62373), .ZN(n27712) );
  INV_X1 U32183 ( .A(n27712), .ZN(p_wishbone_bd_ram_n24120) );
  INV_X1 U32184 ( .A(n62372), .ZN(n27714) );
  INV_X1 U32185 ( .A(n27714), .ZN(p_wishbone_bd_ram_n24118) );
  INV_X1 U32186 ( .A(n62371), .ZN(n27716) );
  INV_X1 U32187 ( .A(n27716), .ZN(p_wishbone_bd_ram_n24115) );
  INV_X1 U32188 ( .A(n62370), .ZN(n27718) );
  INV_X1 U32189 ( .A(n27718), .ZN(p_wishbone_bd_ram_n24113) );
  INV_X1 U32190 ( .A(n62369), .ZN(n27720) );
  INV_X1 U32191 ( .A(n27720), .ZN(p_wishbone_bd_ram_n24112) );
  INV_X1 U32192 ( .A(n62368), .ZN(n27722) );
  INV_X1 U32193 ( .A(n27722), .ZN(p_wishbone_bd_ram_n24111) );
  INV_X1 U32194 ( .A(n62367), .ZN(n27724) );
  INV_X1 U32195 ( .A(n27724), .ZN(p_wishbone_bd_ram_n24110) );
  INV_X1 U32196 ( .A(n62366), .ZN(n27726) );
  INV_X1 U32197 ( .A(n27726), .ZN(p_wishbone_bd_ram_n24109) );
  INV_X1 U32198 ( .A(n62365), .ZN(n27728) );
  INV_X1 U32199 ( .A(n27728), .ZN(p_wishbone_bd_ram_n24108) );
  INV_X1 U32200 ( .A(n62364), .ZN(n27730) );
  INV_X1 U32201 ( .A(n27730), .ZN(p_wishbone_bd_ram_n24107) );
  INV_X1 U32202 ( .A(n62363), .ZN(n27732) );
  INV_X1 U32203 ( .A(n27732), .ZN(p_wishbone_bd_ram_n24106) );
  INV_X1 U32204 ( .A(n62362), .ZN(n27734) );
  INV_X1 U32205 ( .A(n27734), .ZN(p_wishbone_bd_ram_n24105) );
  INV_X1 U32206 ( .A(n62361), .ZN(n27736) );
  INV_X1 U32207 ( .A(n27736), .ZN(p_wishbone_bd_ram_n24104) );
  INV_X1 U32208 ( .A(n62360), .ZN(n27738) );
  INV_X1 U32209 ( .A(n27738), .ZN(p_wishbone_bd_ram_n24102) );
  INV_X1 U32210 ( .A(n62359), .ZN(n27740) );
  INV_X1 U32211 ( .A(n27740), .ZN(p_wishbone_bd_ram_n24099) );
  INV_X1 U32212 ( .A(n62358), .ZN(n27742) );
  INV_X1 U32213 ( .A(n27742), .ZN(p_wishbone_bd_ram_n24097) );
  INV_X1 U32214 ( .A(n62357), .ZN(n27744) );
  INV_X1 U32215 ( .A(n27744), .ZN(p_wishbone_bd_ram_n24096) );
  INV_X1 U32216 ( .A(n62356), .ZN(n27746) );
  INV_X1 U32217 ( .A(n27746), .ZN(p_wishbone_bd_ram_n24095) );
  INV_X1 U32218 ( .A(n62355), .ZN(n27748) );
  INV_X1 U32219 ( .A(n27748), .ZN(p_wishbone_bd_ram_n24094) );
  INV_X1 U32220 ( .A(n62354), .ZN(n27750) );
  INV_X1 U32221 ( .A(n27750), .ZN(p_wishbone_bd_ram_n24093) );
  INV_X1 U32222 ( .A(n62353), .ZN(n27752) );
  INV_X1 U32223 ( .A(n27752), .ZN(p_wishbone_bd_ram_n24092) );
  INV_X1 U32224 ( .A(n62352), .ZN(n27754) );
  INV_X1 U32225 ( .A(n27754), .ZN(p_wishbone_bd_ram_n24091) );
  INV_X1 U32226 ( .A(n62351), .ZN(n27756) );
  INV_X1 U32227 ( .A(n27756), .ZN(p_wishbone_bd_ram_n24090) );
  INV_X1 U32228 ( .A(n62350), .ZN(n27758) );
  INV_X1 U32229 ( .A(n27758), .ZN(p_wishbone_bd_ram_n24089) );
  INV_X1 U32230 ( .A(n62349), .ZN(n27760) );
  INV_X1 U32231 ( .A(n27760), .ZN(p_wishbone_bd_ram_n24087) );
  INV_X1 U32232 ( .A(n62348), .ZN(n27762) );
  INV_X1 U32233 ( .A(n27762), .ZN(p_wishbone_bd_ram_n24085) );
  INV_X1 U32234 ( .A(n62347), .ZN(n27764) );
  INV_X1 U32235 ( .A(n27764), .ZN(p_wishbone_bd_ram_n24084) );
  INV_X1 U32236 ( .A(n62346), .ZN(n27766) );
  INV_X1 U32237 ( .A(n27766), .ZN(p_wishbone_bd_ram_n24082) );
  INV_X1 U32238 ( .A(n62345), .ZN(n27768) );
  INV_X1 U32239 ( .A(n27768), .ZN(p_wishbone_bd_ram_n24080) );
  INV_X1 U32240 ( .A(n62344), .ZN(n27770) );
  INV_X1 U32241 ( .A(n27770), .ZN(p_wishbone_bd_ram_n24078) );
  INV_X1 U32242 ( .A(n62343), .ZN(n27772) );
  INV_X1 U32243 ( .A(n27772), .ZN(p_wishbone_bd_ram_n24075) );
  INV_X1 U32244 ( .A(n62342), .ZN(n27774) );
  INV_X1 U32245 ( .A(n27774), .ZN(p_wishbone_bd_ram_n24073) );
  INV_X1 U32246 ( .A(n62341), .ZN(n27776) );
  INV_X1 U32247 ( .A(n27776), .ZN(p_wishbone_bd_ram_n24072) );
  INV_X1 U32248 ( .A(n62340), .ZN(n27778) );
  INV_X1 U32249 ( .A(n27778), .ZN(p_wishbone_bd_ram_n24070) );
  INV_X1 U32250 ( .A(n62339), .ZN(n27780) );
  INV_X1 U32251 ( .A(n27780), .ZN(p_wishbone_bd_ram_n24067) );
  INV_X1 U32252 ( .A(n62338), .ZN(n27782) );
  INV_X1 U32253 ( .A(n27782), .ZN(p_wishbone_bd_ram_n24065) );
  INV_X1 U32254 ( .A(n62337), .ZN(n27784) );
  INV_X1 U32255 ( .A(n27784), .ZN(p_wishbone_bd_ram_n24064) );
  INV_X1 U32256 ( .A(n62336), .ZN(n27786) );
  INV_X1 U32257 ( .A(n27786), .ZN(p_wishbone_bd_ram_n24062) );
  INV_X1 U32258 ( .A(n62335), .ZN(n27788) );
  INV_X1 U32259 ( .A(n27788), .ZN(p_wishbone_bd_ram_n24059) );
  INV_X1 U32260 ( .A(n62334), .ZN(n27790) );
  INV_X1 U32261 ( .A(n27790), .ZN(p_wishbone_bd_ram_n24057) );
  INV_X1 U32262 ( .A(n62333), .ZN(n27792) );
  INV_X1 U32263 ( .A(n27792), .ZN(p_wishbone_bd_ram_n24055) );
  INV_X1 U32264 ( .A(n62332), .ZN(n27794) );
  INV_X1 U32265 ( .A(n27794), .ZN(p_wishbone_bd_ram_n24053) );
  INV_X1 U32266 ( .A(n62331), .ZN(n27796) );
  INV_X1 U32267 ( .A(n27796), .ZN(p_wishbone_bd_ram_n24052) );
  INV_X1 U32268 ( .A(n62330), .ZN(n27798) );
  INV_X1 U32269 ( .A(n27798), .ZN(p_wishbone_bd_ram_n24050) );
  INV_X1 U32270 ( .A(n62329), .ZN(n27800) );
  INV_X1 U32271 ( .A(n27800), .ZN(p_wishbone_bd_ram_n24048) );
  INV_X1 U32272 ( .A(n62328), .ZN(n27802) );
  INV_X1 U32273 ( .A(n27802), .ZN(p_wishbone_bd_ram_n24047) );
  INV_X1 U32274 ( .A(n62327), .ZN(n27804) );
  INV_X1 U32275 ( .A(n27804), .ZN(p_wishbone_bd_ram_n24046) );
  INV_X1 U32276 ( .A(n62326), .ZN(n27806) );
  INV_X1 U32277 ( .A(n27806), .ZN(p_wishbone_bd_ram_n24045) );
  INV_X1 U32278 ( .A(n62325), .ZN(n27808) );
  INV_X1 U32279 ( .A(n27808), .ZN(p_wishbone_bd_ram_n24044) );
  INV_X1 U32280 ( .A(n62324), .ZN(n27810) );
  INV_X1 U32281 ( .A(n27810), .ZN(p_wishbone_bd_ram_n24043) );
  INV_X1 U32282 ( .A(n62323), .ZN(n27812) );
  INV_X1 U32283 ( .A(n27812), .ZN(p_wishbone_bd_ram_n24042) );
  INV_X1 U32284 ( .A(n62322), .ZN(n27814) );
  INV_X1 U32285 ( .A(n27814), .ZN(p_wishbone_bd_ram_n24041) );
  INV_X1 U32286 ( .A(n62321), .ZN(n27816) );
  INV_X1 U32287 ( .A(n27816), .ZN(p_wishbone_bd_ram_n24040) );
  INV_X1 U32288 ( .A(n62320), .ZN(n27818) );
  INV_X1 U32289 ( .A(n27818), .ZN(p_wishbone_bd_ram_n24039) );
  INV_X1 U32290 ( .A(n62319), .ZN(n27820) );
  INV_X1 U32291 ( .A(n27820), .ZN(p_wishbone_bd_ram_n24038) );
  INV_X1 U32292 ( .A(n62318), .ZN(n27822) );
  INV_X1 U32293 ( .A(n27822), .ZN(p_wishbone_bd_ram_n24037) );
  INV_X1 U32294 ( .A(n62317), .ZN(n27824) );
  INV_X1 U32295 ( .A(n27824), .ZN(p_wishbone_bd_ram_n24036) );
  INV_X1 U32296 ( .A(n62316), .ZN(n27826) );
  INV_X1 U32297 ( .A(n27826), .ZN(p_wishbone_bd_ram_n24035) );
  INV_X1 U32298 ( .A(n62315), .ZN(n27828) );
  INV_X1 U32299 ( .A(n27828), .ZN(p_wishbone_bd_ram_n24034) );
  INV_X1 U32300 ( .A(n62314), .ZN(n27830) );
  INV_X1 U32301 ( .A(n27830), .ZN(p_wishbone_bd_ram_n24033) );
  INV_X1 U32302 ( .A(n62313), .ZN(n27832) );
  INV_X1 U32303 ( .A(n27832), .ZN(p_wishbone_bd_ram_n24032) );
  INV_X1 U32304 ( .A(n62312), .ZN(n27834) );
  INV_X1 U32305 ( .A(n27834), .ZN(p_wishbone_bd_ram_n24031) );
  INV_X1 U32306 ( .A(n62311), .ZN(n27836) );
  INV_X1 U32307 ( .A(n27836), .ZN(p_wishbone_bd_ram_n24030) );
  INV_X1 U32308 ( .A(n62310), .ZN(n27838) );
  INV_X1 U32309 ( .A(n27838), .ZN(p_wishbone_bd_ram_n24029) );
  INV_X1 U32310 ( .A(n62309), .ZN(n27840) );
  INV_X1 U32311 ( .A(n27840), .ZN(p_wishbone_bd_ram_n24028) );
  INV_X1 U32312 ( .A(n62308), .ZN(n27842) );
  INV_X1 U32313 ( .A(n27842), .ZN(p_wishbone_bd_ram_n24027) );
  INV_X1 U32314 ( .A(n62307), .ZN(n27844) );
  INV_X1 U32315 ( .A(n27844), .ZN(p_wishbone_bd_ram_n24026) );
  INV_X1 U32316 ( .A(n62306), .ZN(n27846) );
  INV_X1 U32317 ( .A(n27846), .ZN(p_wishbone_bd_ram_n24025) );
  INV_X1 U32318 ( .A(n62305), .ZN(n27848) );
  INV_X1 U32319 ( .A(n27848), .ZN(p_wishbone_bd_ram_n24023) );
  INV_X1 U32320 ( .A(n62304), .ZN(n27850) );
  INV_X1 U32321 ( .A(n27850), .ZN(p_wishbone_bd_ram_n24021) );
  INV_X1 U32322 ( .A(n62303), .ZN(n27852) );
  INV_X1 U32323 ( .A(n27852), .ZN(p_wishbone_bd_ram_n24020) );
  INV_X1 U32324 ( .A(n62302), .ZN(n27854) );
  INV_X1 U32325 ( .A(n27854), .ZN(p_wishbone_bd_ram_n24018) );
  INV_X1 U32326 ( .A(n62301), .ZN(n27856) );
  INV_X1 U32327 ( .A(n27856), .ZN(p_wishbone_bd_ram_n24016) );
  INV_X1 U32328 ( .A(n62300), .ZN(n27858) );
  INV_X1 U32329 ( .A(n27858), .ZN(p_wishbone_bd_ram_n24015) );
  INV_X1 U32330 ( .A(n62299), .ZN(n27860) );
  INV_X1 U32331 ( .A(n27860), .ZN(p_wishbone_bd_ram_n24014) );
  INV_X1 U32332 ( .A(n62298), .ZN(n27862) );
  INV_X1 U32333 ( .A(n27862), .ZN(p_wishbone_bd_ram_n24013) );
  INV_X1 U32334 ( .A(n62297), .ZN(n27864) );
  INV_X1 U32335 ( .A(n27864), .ZN(p_wishbone_bd_ram_n24012) );
  INV_X1 U32336 ( .A(n62296), .ZN(n27866) );
  INV_X1 U32337 ( .A(n27866), .ZN(p_wishbone_bd_ram_n24011) );
  INV_X1 U32338 ( .A(n62295), .ZN(n27868) );
  INV_X1 U32339 ( .A(n27868), .ZN(p_wishbone_bd_ram_n24010) );
  INV_X1 U32340 ( .A(n62294), .ZN(n27870) );
  INV_X1 U32341 ( .A(n27870), .ZN(p_wishbone_bd_ram_n24009) );
  INV_X1 U32342 ( .A(n62293), .ZN(n27872) );
  INV_X1 U32343 ( .A(n27872), .ZN(p_wishbone_bd_ram_n24008) );
  INV_X1 U32344 ( .A(n62292), .ZN(n27874) );
  INV_X1 U32345 ( .A(n27874), .ZN(p_wishbone_bd_ram_n24007) );
  INV_X1 U32346 ( .A(n62291), .ZN(n27876) );
  INV_X1 U32347 ( .A(n27876), .ZN(p_wishbone_bd_ram_n24006) );
  INV_X1 U32348 ( .A(n62290), .ZN(n27878) );
  INV_X1 U32349 ( .A(n27878), .ZN(p_wishbone_bd_ram_n24005) );
  INV_X1 U32350 ( .A(n62289), .ZN(n27880) );
  INV_X1 U32351 ( .A(n27880), .ZN(p_wishbone_bd_ram_n24004) );
  INV_X1 U32352 ( .A(n62288), .ZN(n27882) );
  INV_X1 U32353 ( .A(n27882), .ZN(p_wishbone_bd_ram_n24003) );
  INV_X1 U32354 ( .A(n62287), .ZN(n27884) );
  INV_X1 U32355 ( .A(n27884), .ZN(p_wishbone_bd_ram_n24002) );
  INV_X1 U32356 ( .A(n62286), .ZN(n27886) );
  INV_X1 U32357 ( .A(n27886), .ZN(p_wishbone_bd_ram_n24001) );
  INV_X1 U32358 ( .A(n62285), .ZN(n27888) );
  INV_X1 U32359 ( .A(n27888), .ZN(p_wishbone_bd_ram_n23999) );
  INV_X1 U32360 ( .A(n62284), .ZN(n27890) );
  INV_X1 U32361 ( .A(n27890), .ZN(p_wishbone_bd_ram_n23997) );
  INV_X1 U32362 ( .A(n62283), .ZN(n27892) );
  INV_X1 U32363 ( .A(n27892), .ZN(p_wishbone_bd_ram_n23996) );
  INV_X1 U32364 ( .A(n62282), .ZN(n27894) );
  INV_X1 U32365 ( .A(n27894), .ZN(p_wishbone_bd_ram_n23994) );
  INV_X1 U32366 ( .A(n62281), .ZN(n27896) );
  INV_X1 U32367 ( .A(n27896), .ZN(p_wishbone_bd_ram_n23991) );
  INV_X1 U32368 ( .A(n62280), .ZN(n27898) );
  INV_X1 U32369 ( .A(n27898), .ZN(p_wishbone_bd_ram_n23989) );
  INV_X1 U32370 ( .A(n62279), .ZN(n27900) );
  INV_X1 U32371 ( .A(n27900), .ZN(p_wishbone_bd_ram_n23988) );
  INV_X1 U32372 ( .A(n62278), .ZN(n27902) );
  INV_X1 U32373 ( .A(n27902), .ZN(p_wishbone_bd_ram_n23986) );
  INV_X1 U32374 ( .A(n62277), .ZN(n27904) );
  INV_X1 U32375 ( .A(n27904), .ZN(p_wishbone_bd_ram_n23984) );
  INV_X1 U32376 ( .A(n62276), .ZN(n27906) );
  INV_X1 U32377 ( .A(n27906), .ZN(p_wishbone_bd_ram_n23983) );
  INV_X1 U32378 ( .A(n62275), .ZN(n27908) );
  INV_X1 U32379 ( .A(n27908), .ZN(p_wishbone_bd_ram_n23982) );
  INV_X1 U32380 ( .A(n62274), .ZN(n27910) );
  INV_X1 U32381 ( .A(n27910), .ZN(p_wishbone_bd_ram_n23981) );
  INV_X1 U32382 ( .A(n62273), .ZN(n27912) );
  INV_X1 U32383 ( .A(n27912), .ZN(p_wishbone_bd_ram_n23980) );
  INV_X1 U32384 ( .A(n62272), .ZN(n27914) );
  INV_X1 U32385 ( .A(n27914), .ZN(p_wishbone_bd_ram_n23979) );
  INV_X1 U32386 ( .A(n62271), .ZN(n27916) );
  INV_X1 U32387 ( .A(n27916), .ZN(p_wishbone_bd_ram_n23978) );
  INV_X1 U32388 ( .A(n62270), .ZN(n27918) );
  INV_X1 U32389 ( .A(n27918), .ZN(p_wishbone_bd_ram_n23977) );
  INV_X1 U32390 ( .A(n62269), .ZN(n27920) );
  INV_X1 U32391 ( .A(n27920), .ZN(p_wishbone_bd_ram_n23976) );
  INV_X1 U32392 ( .A(n62268), .ZN(n27922) );
  INV_X1 U32393 ( .A(n27922), .ZN(p_wishbone_bd_ram_n23975) );
  INV_X1 U32394 ( .A(n62267), .ZN(n27924) );
  INV_X1 U32395 ( .A(n27924), .ZN(p_wishbone_bd_ram_n23974) );
  INV_X1 U32396 ( .A(n62266), .ZN(n27926) );
  INV_X1 U32397 ( .A(n27926), .ZN(p_wishbone_bd_ram_n23973) );
  INV_X1 U32398 ( .A(n62265), .ZN(n27928) );
  INV_X1 U32399 ( .A(n27928), .ZN(p_wishbone_bd_ram_n23972) );
  INV_X1 U32400 ( .A(n62264), .ZN(n27930) );
  INV_X1 U32401 ( .A(n27930), .ZN(p_wishbone_bd_ram_n23971) );
  INV_X1 U32402 ( .A(n62263), .ZN(n27932) );
  INV_X1 U32403 ( .A(n27932), .ZN(p_wishbone_bd_ram_n23970) );
  INV_X1 U32404 ( .A(n62262), .ZN(n27934) );
  INV_X1 U32405 ( .A(n27934), .ZN(p_wishbone_bd_ram_n23969) );
  INV_X1 U32406 ( .A(n62261), .ZN(n27936) );
  INV_X1 U32407 ( .A(n27936), .ZN(p_wishbone_bd_ram_n23968) );
  INV_X1 U32408 ( .A(n62260), .ZN(n27938) );
  INV_X1 U32409 ( .A(n27938), .ZN(p_wishbone_bd_ram_n23967) );
  INV_X1 U32410 ( .A(n62259), .ZN(n27940) );
  INV_X1 U32411 ( .A(n27940), .ZN(p_wishbone_bd_ram_n23966) );
  INV_X1 U32412 ( .A(n62258), .ZN(n27942) );
  INV_X1 U32413 ( .A(n27942), .ZN(p_wishbone_bd_ram_n23965) );
  INV_X1 U32414 ( .A(n62257), .ZN(n27944) );
  INV_X1 U32415 ( .A(n27944), .ZN(p_wishbone_bd_ram_n23964) );
  INV_X1 U32416 ( .A(n62256), .ZN(n27946) );
  INV_X1 U32417 ( .A(n27946), .ZN(p_wishbone_bd_ram_n23963) );
  INV_X1 U32418 ( .A(n62255), .ZN(n27948) );
  INV_X1 U32419 ( .A(n27948), .ZN(p_wishbone_bd_ram_n23962) );
  INV_X1 U32420 ( .A(n62254), .ZN(n27950) );
  INV_X1 U32421 ( .A(n27950), .ZN(p_wishbone_bd_ram_n23961) );
  INV_X1 U32422 ( .A(n62253), .ZN(n27952) );
  INV_X1 U32423 ( .A(n27952), .ZN(p_wishbone_bd_ram_n23960) );
  INV_X1 U32424 ( .A(n62252), .ZN(n27954) );
  INV_X1 U32425 ( .A(n27954), .ZN(p_wishbone_bd_ram_n23959) );
  INV_X1 U32426 ( .A(n62251), .ZN(n27956) );
  INV_X1 U32427 ( .A(n27956), .ZN(p_wishbone_bd_ram_n23958) );
  INV_X1 U32428 ( .A(n62250), .ZN(n27958) );
  INV_X1 U32429 ( .A(n27958), .ZN(p_wishbone_bd_ram_n23957) );
  INV_X1 U32430 ( .A(n62249), .ZN(n27960) );
  INV_X1 U32431 ( .A(n27960), .ZN(p_wishbone_bd_ram_n23956) );
  INV_X1 U32432 ( .A(n62248), .ZN(n27962) );
  INV_X1 U32433 ( .A(n27962), .ZN(p_wishbone_bd_ram_n23955) );
  INV_X1 U32434 ( .A(n62247), .ZN(n27964) );
  INV_X1 U32435 ( .A(n27964), .ZN(p_wishbone_bd_ram_n23954) );
  INV_X1 U32436 ( .A(n62246), .ZN(n27966) );
  INV_X1 U32437 ( .A(n27966), .ZN(p_wishbone_bd_ram_n23953) );
  INV_X1 U32438 ( .A(n62245), .ZN(n27968) );
  INV_X1 U32439 ( .A(n27968), .ZN(p_wishbone_bd_ram_n23952) );
  INV_X1 U32440 ( .A(n62244), .ZN(n27970) );
  INV_X1 U32441 ( .A(n27970), .ZN(p_wishbone_bd_ram_n23951) );
  INV_X1 U32442 ( .A(n62243), .ZN(n27972) );
  INV_X1 U32443 ( .A(n27972), .ZN(p_wishbone_bd_ram_n23950) );
  INV_X1 U32444 ( .A(n62242), .ZN(n27974) );
  INV_X1 U32445 ( .A(n27974), .ZN(p_wishbone_bd_ram_n23949) );
  INV_X1 U32446 ( .A(n62241), .ZN(n27976) );
  INV_X1 U32447 ( .A(n27976), .ZN(p_wishbone_bd_ram_n23948) );
  INV_X1 U32448 ( .A(n62240), .ZN(n27978) );
  INV_X1 U32449 ( .A(n27978), .ZN(p_wishbone_bd_ram_n23947) );
  INV_X1 U32450 ( .A(n62239), .ZN(n27980) );
  INV_X1 U32451 ( .A(n27980), .ZN(p_wishbone_bd_ram_n23946) );
  INV_X1 U32452 ( .A(n62238), .ZN(n27982) );
  INV_X1 U32453 ( .A(n27982), .ZN(p_wishbone_bd_ram_n23945) );
  INV_X1 U32454 ( .A(n62237), .ZN(n27984) );
  INV_X1 U32455 ( .A(n27984), .ZN(p_wishbone_bd_ram_n23944) );
  INV_X1 U32456 ( .A(n62236), .ZN(n27986) );
  INV_X1 U32457 ( .A(n27986), .ZN(p_wishbone_bd_ram_n23943) );
  INV_X1 U32458 ( .A(n62235), .ZN(n27988) );
  INV_X1 U32459 ( .A(n27988), .ZN(p_wishbone_bd_ram_n23942) );
  INV_X1 U32460 ( .A(n62234), .ZN(n27990) );
  INV_X1 U32461 ( .A(n27990), .ZN(p_wishbone_bd_ram_n23941) );
  INV_X1 U32462 ( .A(n62233), .ZN(n27992) );
  INV_X1 U32463 ( .A(n27992), .ZN(p_wishbone_bd_ram_n23940) );
  INV_X1 U32464 ( .A(n62232), .ZN(n27994) );
  INV_X1 U32465 ( .A(n27994), .ZN(p_wishbone_bd_ram_n23939) );
  INV_X1 U32466 ( .A(n62231), .ZN(n27996) );
  INV_X1 U32467 ( .A(n27996), .ZN(p_wishbone_bd_ram_n23938) );
  INV_X1 U32468 ( .A(n62230), .ZN(n27998) );
  INV_X1 U32469 ( .A(n27998), .ZN(p_wishbone_bd_ram_n23937) );
  INV_X1 U32470 ( .A(n62229), .ZN(n28000) );
  INV_X1 U32471 ( .A(n28000), .ZN(p_wishbone_bd_ram_n23936) );
  INV_X1 U32472 ( .A(n62228), .ZN(n28002) );
  INV_X1 U32473 ( .A(n28002), .ZN(p_wishbone_bd_ram_n23935) );
  INV_X1 U32474 ( .A(n62227), .ZN(n28004) );
  INV_X1 U32475 ( .A(n28004), .ZN(p_wishbone_bd_ram_n23934) );
  INV_X1 U32476 ( .A(n62226), .ZN(n28006) );
  INV_X1 U32477 ( .A(n28006), .ZN(p_wishbone_bd_ram_n23933) );
  INV_X1 U32478 ( .A(n62225), .ZN(n28008) );
  INV_X1 U32479 ( .A(n28008), .ZN(p_wishbone_bd_ram_n23932) );
  INV_X1 U32480 ( .A(n62224), .ZN(n28010) );
  INV_X1 U32481 ( .A(n28010), .ZN(p_wishbone_bd_ram_n23931) );
  INV_X1 U32482 ( .A(n62223), .ZN(n28012) );
  INV_X1 U32483 ( .A(n28012), .ZN(p_wishbone_bd_ram_n23930) );
  INV_X1 U32484 ( .A(n62222), .ZN(n28014) );
  INV_X1 U32485 ( .A(n28014), .ZN(p_wishbone_bd_ram_n23929) );
  INV_X1 U32486 ( .A(n62221), .ZN(n28016) );
  INV_X1 U32487 ( .A(n28016), .ZN(p_wishbone_bd_ram_n23928) );
  INV_X1 U32488 ( .A(n62220), .ZN(n28018) );
  INV_X1 U32489 ( .A(n28018), .ZN(p_wishbone_bd_ram_n23927) );
  INV_X1 U32490 ( .A(n62219), .ZN(n28020) );
  INV_X1 U32491 ( .A(n28020), .ZN(p_wishbone_bd_ram_n23926) );
  INV_X1 U32492 ( .A(n62218), .ZN(n28022) );
  INV_X1 U32493 ( .A(n28022), .ZN(p_wishbone_bd_ram_n23925) );
  INV_X1 U32494 ( .A(n62217), .ZN(n28024) );
  INV_X1 U32495 ( .A(n28024), .ZN(p_wishbone_bd_ram_n23924) );
  INV_X1 U32496 ( .A(n62216), .ZN(n28026) );
  INV_X1 U32497 ( .A(n28026), .ZN(p_wishbone_bd_ram_n23923) );
  INV_X1 U32498 ( .A(n62215), .ZN(n28028) );
  INV_X1 U32499 ( .A(n28028), .ZN(p_wishbone_bd_ram_n23922) );
  INV_X1 U32500 ( .A(n62214), .ZN(n28030) );
  INV_X1 U32501 ( .A(n28030), .ZN(p_wishbone_bd_ram_n23921) );
  INV_X1 U32502 ( .A(n62213), .ZN(n28032) );
  INV_X1 U32503 ( .A(n28032), .ZN(p_wishbone_bd_ram_n23920) );
  INV_X1 U32504 ( .A(n62212), .ZN(n28034) );
  INV_X1 U32505 ( .A(n28034), .ZN(p_wishbone_bd_ram_n23919) );
  INV_X1 U32506 ( .A(n62211), .ZN(n28036) );
  INV_X1 U32507 ( .A(n28036), .ZN(p_wishbone_bd_ram_n23918) );
  INV_X1 U32508 ( .A(n62210), .ZN(n28038) );
  INV_X1 U32509 ( .A(n28038), .ZN(p_wishbone_bd_ram_n23917) );
  INV_X1 U32510 ( .A(n62209), .ZN(n28040) );
  INV_X1 U32511 ( .A(n28040), .ZN(p_wishbone_bd_ram_n23916) );
  INV_X1 U32512 ( .A(n62208), .ZN(n28042) );
  INV_X1 U32513 ( .A(n28042), .ZN(p_wishbone_bd_ram_n23915) );
  INV_X1 U32514 ( .A(n62207), .ZN(n28044) );
  INV_X1 U32515 ( .A(n28044), .ZN(p_wishbone_bd_ram_n23914) );
  INV_X1 U32516 ( .A(n62206), .ZN(n28046) );
  INV_X1 U32517 ( .A(n28046), .ZN(p_wishbone_bd_ram_n23913) );
  INV_X1 U32518 ( .A(n62205), .ZN(n28048) );
  INV_X1 U32519 ( .A(n28048), .ZN(p_wishbone_bd_ram_n23912) );
  INV_X1 U32520 ( .A(n62204), .ZN(n28050) );
  INV_X1 U32521 ( .A(n28050), .ZN(p_wishbone_bd_ram_n23911) );
  INV_X1 U32522 ( .A(n62203), .ZN(n28052) );
  INV_X1 U32523 ( .A(n28052), .ZN(p_wishbone_bd_ram_n23910) );
  INV_X1 U32524 ( .A(n62202), .ZN(n28054) );
  INV_X1 U32525 ( .A(n28054), .ZN(p_wishbone_bd_ram_n23909) );
  INV_X1 U32526 ( .A(n62201), .ZN(n28056) );
  INV_X1 U32527 ( .A(n28056), .ZN(p_wishbone_bd_ram_n23908) );
  INV_X1 U32528 ( .A(n62200), .ZN(n28058) );
  INV_X1 U32529 ( .A(n28058), .ZN(p_wishbone_bd_ram_n23907) );
  INV_X1 U32530 ( .A(n62199), .ZN(n28060) );
  INV_X1 U32531 ( .A(n28060), .ZN(p_wishbone_bd_ram_n23906) );
  INV_X1 U32532 ( .A(n62198), .ZN(n28062) );
  INV_X1 U32533 ( .A(n28062), .ZN(p_wishbone_bd_ram_n23905) );
  INV_X1 U32534 ( .A(n62197), .ZN(n28064) );
  INV_X1 U32535 ( .A(n28064), .ZN(p_wishbone_bd_ram_n23904) );
  INV_X1 U32536 ( .A(n62196), .ZN(n28066) );
  INV_X1 U32537 ( .A(n28066), .ZN(p_wishbone_bd_ram_n23903) );
  INV_X1 U32538 ( .A(n62195), .ZN(n28068) );
  INV_X1 U32539 ( .A(n28068), .ZN(p_wishbone_bd_ram_n23902) );
  INV_X1 U32540 ( .A(n62194), .ZN(n28070) );
  INV_X1 U32541 ( .A(n28070), .ZN(p_wishbone_bd_ram_n23901) );
  INV_X1 U32542 ( .A(n62193), .ZN(n28072) );
  INV_X1 U32543 ( .A(n28072), .ZN(p_wishbone_bd_ram_n23900) );
  INV_X1 U32544 ( .A(n62192), .ZN(n28074) );
  INV_X1 U32545 ( .A(n28074), .ZN(p_wishbone_bd_ram_n23899) );
  INV_X1 U32546 ( .A(n62191), .ZN(n28076) );
  INV_X1 U32547 ( .A(n28076), .ZN(p_wishbone_bd_ram_n23898) );
  INV_X1 U32548 ( .A(n62190), .ZN(n28078) );
  INV_X1 U32549 ( .A(n28078), .ZN(p_wishbone_bd_ram_n23897) );
  INV_X1 U32550 ( .A(n62189), .ZN(n28080) );
  INV_X1 U32551 ( .A(n28080), .ZN(p_wishbone_bd_ram_n23896) );
  INV_X1 U32552 ( .A(n62188), .ZN(n28082) );
  INV_X1 U32553 ( .A(n28082), .ZN(p_wishbone_bd_ram_n23895) );
  INV_X1 U32554 ( .A(n62187), .ZN(n28084) );
  INV_X1 U32555 ( .A(n28084), .ZN(p_wishbone_bd_ram_n23894) );
  INV_X1 U32556 ( .A(n62186), .ZN(n28086) );
  INV_X1 U32557 ( .A(n28086), .ZN(p_wishbone_bd_ram_n23893) );
  INV_X1 U32558 ( .A(n62185), .ZN(n28088) );
  INV_X1 U32559 ( .A(n28088), .ZN(p_wishbone_bd_ram_n23892) );
  INV_X1 U32560 ( .A(n62184), .ZN(n28090) );
  INV_X1 U32561 ( .A(n28090), .ZN(p_wishbone_bd_ram_n23891) );
  INV_X1 U32562 ( .A(n62183), .ZN(n28092) );
  INV_X1 U32563 ( .A(n28092), .ZN(p_wishbone_bd_ram_n23890) );
  INV_X1 U32564 ( .A(n62182), .ZN(n28094) );
  INV_X1 U32565 ( .A(n28094), .ZN(p_wishbone_bd_ram_n23889) );
  INV_X1 U32566 ( .A(n62181), .ZN(n28096) );
  INV_X1 U32567 ( .A(n28096), .ZN(p_wishbone_bd_ram_n23888) );
  INV_X1 U32568 ( .A(n62180), .ZN(n28098) );
  INV_X1 U32569 ( .A(n28098), .ZN(p_wishbone_bd_ram_n23887) );
  INV_X1 U32570 ( .A(n62179), .ZN(n28100) );
  INV_X1 U32571 ( .A(n28100), .ZN(p_wishbone_bd_ram_n23886) );
  INV_X1 U32572 ( .A(n62178), .ZN(n28102) );
  INV_X1 U32573 ( .A(n28102), .ZN(p_wishbone_bd_ram_n23885) );
  INV_X1 U32574 ( .A(n62177), .ZN(n28104) );
  INV_X1 U32575 ( .A(n28104), .ZN(p_wishbone_bd_ram_n23884) );
  INV_X1 U32576 ( .A(n62176), .ZN(n28106) );
  INV_X1 U32577 ( .A(n28106), .ZN(p_wishbone_bd_ram_n23883) );
  INV_X1 U32578 ( .A(n62175), .ZN(n28108) );
  INV_X1 U32579 ( .A(n28108), .ZN(p_wishbone_bd_ram_n23882) );
  INV_X1 U32580 ( .A(n62174), .ZN(n28110) );
  INV_X1 U32581 ( .A(n28110), .ZN(p_wishbone_bd_ram_n23881) );
  INV_X1 U32582 ( .A(n62173), .ZN(n28112) );
  INV_X1 U32583 ( .A(n28112), .ZN(p_wishbone_bd_ram_n23880) );
  INV_X1 U32584 ( .A(n62172), .ZN(n28114) );
  INV_X1 U32585 ( .A(n28114), .ZN(p_wishbone_bd_ram_n23879) );
  INV_X1 U32586 ( .A(n62171), .ZN(n28116) );
  INV_X1 U32587 ( .A(n28116), .ZN(p_wishbone_bd_ram_n23878) );
  INV_X1 U32588 ( .A(n62170), .ZN(n28118) );
  INV_X1 U32589 ( .A(n28118), .ZN(p_wishbone_bd_ram_n23877) );
  INV_X1 U32590 ( .A(n62169), .ZN(n28120) );
  INV_X1 U32591 ( .A(n28120), .ZN(p_wishbone_bd_ram_n23876) );
  INV_X1 U32592 ( .A(n62168), .ZN(n28122) );
  INV_X1 U32593 ( .A(n28122), .ZN(p_wishbone_bd_ram_n23875) );
  INV_X1 U32594 ( .A(n62167), .ZN(n28124) );
  INV_X1 U32595 ( .A(n28124), .ZN(p_wishbone_bd_ram_n23874) );
  INV_X1 U32596 ( .A(n62166), .ZN(n28126) );
  INV_X1 U32597 ( .A(n28126), .ZN(p_wishbone_bd_ram_n23873) );
  INV_X1 U32598 ( .A(n62165), .ZN(n28128) );
  INV_X1 U32599 ( .A(n28128), .ZN(p_wishbone_bd_ram_n23872) );
  INV_X1 U32600 ( .A(n62164), .ZN(n28130) );
  INV_X1 U32601 ( .A(n28130), .ZN(p_wishbone_bd_ram_n23871) );
  INV_X1 U32602 ( .A(n62163), .ZN(n28132) );
  INV_X1 U32603 ( .A(n28132), .ZN(p_wishbone_bd_ram_n23870) );
  INV_X1 U32604 ( .A(n62162), .ZN(n28134) );
  INV_X1 U32605 ( .A(n28134), .ZN(p_wishbone_bd_ram_n23869) );
  INV_X1 U32606 ( .A(n62161), .ZN(n28136) );
  INV_X1 U32607 ( .A(n28136), .ZN(p_wishbone_bd_ram_n23868) );
  INV_X1 U32608 ( .A(n62160), .ZN(n28138) );
  INV_X1 U32609 ( .A(n28138), .ZN(p_wishbone_bd_ram_n23867) );
  INV_X1 U32610 ( .A(n62159), .ZN(n28140) );
  INV_X1 U32611 ( .A(n28140), .ZN(p_wishbone_bd_ram_n23866) );
  INV_X1 U32612 ( .A(n62158), .ZN(n28142) );
  INV_X1 U32613 ( .A(n28142), .ZN(p_wishbone_bd_ram_n23865) );
  INV_X1 U32614 ( .A(n62157), .ZN(n28144) );
  INV_X1 U32615 ( .A(n28144), .ZN(p_wishbone_bd_ram_n23864) );
  INV_X1 U32616 ( .A(n62156), .ZN(n28146) );
  INV_X1 U32617 ( .A(n28146), .ZN(p_wishbone_bd_ram_n23863) );
  INV_X1 U32618 ( .A(n62155), .ZN(n28148) );
  INV_X1 U32619 ( .A(n28148), .ZN(p_wishbone_bd_ram_n23862) );
  INV_X1 U32620 ( .A(n62154), .ZN(n28150) );
  INV_X1 U32621 ( .A(n28150), .ZN(p_wishbone_bd_ram_n23861) );
  INV_X1 U32622 ( .A(n62153), .ZN(n28152) );
  INV_X1 U32623 ( .A(n28152), .ZN(p_wishbone_bd_ram_n23860) );
  INV_X1 U32624 ( .A(n62152), .ZN(n28154) );
  INV_X1 U32625 ( .A(n28154), .ZN(p_wishbone_bd_ram_n23859) );
  INV_X1 U32626 ( .A(n62151), .ZN(n28156) );
  INV_X1 U32627 ( .A(n28156), .ZN(p_wishbone_bd_ram_n23858) );
  INV_X1 U32628 ( .A(n62150), .ZN(n28158) );
  INV_X1 U32629 ( .A(n28158), .ZN(p_wishbone_bd_ram_n23857) );
  INV_X1 U32630 ( .A(n62149), .ZN(n28160) );
  INV_X1 U32631 ( .A(n28160), .ZN(p_wishbone_bd_ram_n23856) );
  INV_X1 U32632 ( .A(n62148), .ZN(n28162) );
  INV_X1 U32633 ( .A(n28162), .ZN(p_wishbone_bd_ram_n23855) );
  INV_X1 U32634 ( .A(n62147), .ZN(n28164) );
  INV_X1 U32635 ( .A(n28164), .ZN(p_wishbone_bd_ram_n23854) );
  INV_X1 U32636 ( .A(n62146), .ZN(n28166) );
  INV_X1 U32637 ( .A(n28166), .ZN(p_wishbone_bd_ram_n23853) );
  INV_X1 U32638 ( .A(n62145), .ZN(n28168) );
  INV_X1 U32639 ( .A(n28168), .ZN(p_wishbone_bd_ram_n23852) );
  INV_X1 U32640 ( .A(n62144), .ZN(n28170) );
  INV_X1 U32641 ( .A(n28170), .ZN(p_wishbone_bd_ram_n23851) );
  INV_X1 U32642 ( .A(n62143), .ZN(n28172) );
  INV_X1 U32643 ( .A(n28172), .ZN(p_wishbone_bd_ram_n23850) );
  INV_X1 U32644 ( .A(n62142), .ZN(n28174) );
  INV_X1 U32645 ( .A(n28174), .ZN(p_wishbone_bd_ram_n23849) );
  INV_X1 U32646 ( .A(n62141), .ZN(n28176) );
  INV_X1 U32647 ( .A(n28176), .ZN(p_wishbone_bd_ram_n23848) );
  INV_X1 U32648 ( .A(n62140), .ZN(n28178) );
  INV_X1 U32649 ( .A(n28178), .ZN(p_wishbone_bd_ram_n23847) );
  INV_X1 U32650 ( .A(n62139), .ZN(n28180) );
  INV_X1 U32651 ( .A(n28180), .ZN(p_wishbone_bd_ram_n23846) );
  INV_X1 U32652 ( .A(n62138), .ZN(n28182) );
  INV_X1 U32653 ( .A(n28182), .ZN(p_wishbone_bd_ram_n23845) );
  INV_X1 U32654 ( .A(n62137), .ZN(n28184) );
  INV_X1 U32655 ( .A(n28184), .ZN(p_wishbone_bd_ram_n23844) );
  INV_X1 U32656 ( .A(n62136), .ZN(n28186) );
  INV_X1 U32657 ( .A(n28186), .ZN(p_wishbone_bd_ram_n23843) );
  INV_X1 U32658 ( .A(n62135), .ZN(n28188) );
  INV_X1 U32659 ( .A(n28188), .ZN(p_wishbone_bd_ram_n23842) );
  INV_X1 U32660 ( .A(n62134), .ZN(n28190) );
  INV_X1 U32661 ( .A(n28190), .ZN(p_wishbone_bd_ram_n23841) );
  INV_X1 U32662 ( .A(n62133), .ZN(n28192) );
  INV_X1 U32663 ( .A(n28192), .ZN(p_wishbone_bd_ram_n23840) );
  INV_X1 U32664 ( .A(n62132), .ZN(n28194) );
  INV_X1 U32665 ( .A(n28194), .ZN(p_wishbone_bd_ram_n23839) );
  INV_X1 U32666 ( .A(n62131), .ZN(n28196) );
  INV_X1 U32667 ( .A(n28196), .ZN(p_wishbone_bd_ram_n23838) );
  INV_X1 U32668 ( .A(n62130), .ZN(n28198) );
  INV_X1 U32669 ( .A(n28198), .ZN(p_wishbone_bd_ram_n23837) );
  INV_X1 U32670 ( .A(n62129), .ZN(n28200) );
  INV_X1 U32671 ( .A(n28200), .ZN(p_wishbone_bd_ram_n23836) );
  INV_X1 U32672 ( .A(n62128), .ZN(n28202) );
  INV_X1 U32673 ( .A(n28202), .ZN(p_wishbone_bd_ram_n23835) );
  INV_X1 U32674 ( .A(n62127), .ZN(n28204) );
  INV_X1 U32675 ( .A(n28204), .ZN(p_wishbone_bd_ram_n23834) );
  INV_X1 U32676 ( .A(n62126), .ZN(n28206) );
  INV_X1 U32677 ( .A(n28206), .ZN(p_wishbone_bd_ram_n23833) );
  INV_X1 U32678 ( .A(n62125), .ZN(n28208) );
  INV_X1 U32679 ( .A(n28208), .ZN(p_wishbone_bd_ram_n23832) );
  INV_X1 U32680 ( .A(n62124), .ZN(n28210) );
  INV_X1 U32681 ( .A(n28210), .ZN(p_wishbone_bd_ram_n23831) );
  INV_X1 U32682 ( .A(n62123), .ZN(n28212) );
  INV_X1 U32683 ( .A(n28212), .ZN(p_wishbone_bd_ram_n23830) );
  INV_X1 U32684 ( .A(n62122), .ZN(n28214) );
  INV_X1 U32685 ( .A(n28214), .ZN(p_wishbone_bd_ram_n23829) );
  INV_X1 U32686 ( .A(n62121), .ZN(n28216) );
  INV_X1 U32687 ( .A(n28216), .ZN(p_wishbone_bd_ram_n23828) );
  INV_X1 U32688 ( .A(n62120), .ZN(n28218) );
  INV_X1 U32689 ( .A(n28218), .ZN(p_wishbone_bd_ram_n23827) );
  INV_X1 U32690 ( .A(n62119), .ZN(n28220) );
  INV_X1 U32691 ( .A(n28220), .ZN(p_wishbone_bd_ram_n23826) );
  INV_X1 U32692 ( .A(n62118), .ZN(n28222) );
  INV_X1 U32693 ( .A(n28222), .ZN(p_wishbone_bd_ram_n23825) );
  INV_X1 U32694 ( .A(n62117), .ZN(n28224) );
  INV_X1 U32695 ( .A(n28224), .ZN(p_wishbone_bd_ram_n23824) );
  INV_X1 U32696 ( .A(n62116), .ZN(n28226) );
  INV_X1 U32697 ( .A(n28226), .ZN(p_wishbone_bd_ram_n23823) );
  INV_X1 U32698 ( .A(n62115), .ZN(n28228) );
  INV_X1 U32699 ( .A(n28228), .ZN(p_wishbone_bd_ram_n23822) );
  INV_X1 U32700 ( .A(n62114), .ZN(n28230) );
  INV_X1 U32701 ( .A(n28230), .ZN(p_wishbone_bd_ram_n23821) );
  INV_X1 U32702 ( .A(n62113), .ZN(n28232) );
  INV_X1 U32703 ( .A(n28232), .ZN(p_wishbone_bd_ram_n23820) );
  INV_X1 U32704 ( .A(n62112), .ZN(n28234) );
  INV_X1 U32705 ( .A(n28234), .ZN(p_wishbone_bd_ram_n23819) );
  INV_X1 U32706 ( .A(n62111), .ZN(n28236) );
  INV_X1 U32707 ( .A(n28236), .ZN(p_wishbone_bd_ram_n23818) );
  INV_X1 U32708 ( .A(n62110), .ZN(n28238) );
  INV_X1 U32709 ( .A(n28238), .ZN(p_wishbone_bd_ram_n23817) );
  INV_X1 U32710 ( .A(n62109), .ZN(n28240) );
  INV_X1 U32711 ( .A(n28240), .ZN(p_wishbone_bd_ram_n23816) );
  INV_X1 U32712 ( .A(n62108), .ZN(n28242) );
  INV_X1 U32713 ( .A(n28242), .ZN(p_wishbone_bd_ram_n23815) );
  INV_X1 U32714 ( .A(n62107), .ZN(n28244) );
  INV_X1 U32715 ( .A(n28244), .ZN(p_wishbone_bd_ram_n23814) );
  INV_X1 U32716 ( .A(n62106), .ZN(n28246) );
  INV_X1 U32717 ( .A(n28246), .ZN(p_wishbone_bd_ram_n23813) );
  INV_X1 U32718 ( .A(n62105), .ZN(n28248) );
  INV_X1 U32719 ( .A(n28248), .ZN(p_wishbone_bd_ram_n23812) );
  INV_X1 U32720 ( .A(n62104), .ZN(n28250) );
  INV_X1 U32721 ( .A(n28250), .ZN(p_wishbone_bd_ram_n23811) );
  INV_X1 U32722 ( .A(n62103), .ZN(n28252) );
  INV_X1 U32723 ( .A(n28252), .ZN(p_wishbone_bd_ram_n23810) );
  INV_X1 U32724 ( .A(n62102), .ZN(n28254) );
  INV_X1 U32725 ( .A(n28254), .ZN(p_wishbone_bd_ram_n23809) );
  INV_X1 U32726 ( .A(n62101), .ZN(n28256) );
  INV_X1 U32727 ( .A(n28256), .ZN(p_wishbone_bd_ram_n23808) );
  INV_X1 U32728 ( .A(n62100), .ZN(n28258) );
  INV_X1 U32729 ( .A(n28258), .ZN(p_wishbone_bd_ram_n23807) );
  INV_X1 U32730 ( .A(n62099), .ZN(n28260) );
  INV_X1 U32731 ( .A(n28260), .ZN(p_wishbone_bd_ram_n23806) );
  INV_X1 U32732 ( .A(n62098), .ZN(n28262) );
  INV_X1 U32733 ( .A(n28262), .ZN(p_wishbone_bd_ram_n23805) );
  INV_X1 U32734 ( .A(n62097), .ZN(n28264) );
  INV_X1 U32735 ( .A(n28264), .ZN(p_wishbone_bd_ram_n23804) );
  INV_X1 U32736 ( .A(n62096), .ZN(n28266) );
  INV_X1 U32737 ( .A(n28266), .ZN(p_wishbone_bd_ram_n23803) );
  INV_X1 U32738 ( .A(n62095), .ZN(n28268) );
  INV_X1 U32739 ( .A(n28268), .ZN(p_wishbone_bd_ram_n23802) );
  INV_X1 U32740 ( .A(n62094), .ZN(n28270) );
  INV_X1 U32741 ( .A(n28270), .ZN(p_wishbone_bd_ram_n23801) );
  INV_X1 U32742 ( .A(n62093), .ZN(n28272) );
  INV_X1 U32743 ( .A(n28272), .ZN(p_wishbone_bd_ram_n23800) );
  INV_X1 U32744 ( .A(n62092), .ZN(n28274) );
  INV_X1 U32745 ( .A(n28274), .ZN(p_wishbone_bd_ram_n23799) );
  INV_X1 U32746 ( .A(n62091), .ZN(n28276) );
  INV_X1 U32747 ( .A(n28276), .ZN(p_wishbone_bd_ram_n23798) );
  INV_X1 U32748 ( .A(n62090), .ZN(n28278) );
  INV_X1 U32749 ( .A(n28278), .ZN(p_wishbone_bd_ram_n23797) );
  INV_X1 U32750 ( .A(n62089), .ZN(n28280) );
  INV_X1 U32751 ( .A(n28280), .ZN(p_wishbone_bd_ram_n23796) );
  INV_X1 U32752 ( .A(n62088), .ZN(n28282) );
  INV_X1 U32753 ( .A(n28282), .ZN(p_wishbone_bd_ram_n23795) );
  INV_X1 U32754 ( .A(n62087), .ZN(n28284) );
  INV_X1 U32755 ( .A(n28284), .ZN(p_wishbone_bd_ram_n23794) );
  INV_X1 U32756 ( .A(n62086), .ZN(n28286) );
  INV_X1 U32757 ( .A(n28286), .ZN(p_wishbone_bd_ram_n23793) );
  INV_X1 U32758 ( .A(n62085), .ZN(n28288) );
  INV_X1 U32759 ( .A(n28288), .ZN(p_wishbone_bd_ram_n23792) );
  INV_X1 U32760 ( .A(n62084), .ZN(n28290) );
  INV_X1 U32761 ( .A(n28290), .ZN(p_wishbone_bd_ram_n23791) );
  INV_X1 U32762 ( .A(n62083), .ZN(n28292) );
  INV_X1 U32763 ( .A(n28292), .ZN(p_wishbone_bd_ram_n23790) );
  INV_X1 U32764 ( .A(n62082), .ZN(n28294) );
  INV_X1 U32765 ( .A(n28294), .ZN(p_wishbone_bd_ram_n23789) );
  INV_X1 U32766 ( .A(n62081), .ZN(n28296) );
  INV_X1 U32767 ( .A(n28296), .ZN(p_wishbone_bd_ram_n23788) );
  INV_X1 U32768 ( .A(n62080), .ZN(n28298) );
  INV_X1 U32769 ( .A(n28298), .ZN(p_wishbone_bd_ram_n23787) );
  INV_X1 U32770 ( .A(n62079), .ZN(n28300) );
  INV_X1 U32771 ( .A(n28300), .ZN(p_wishbone_bd_ram_n23786) );
  INV_X1 U32772 ( .A(n62078), .ZN(n28302) );
  INV_X1 U32773 ( .A(n28302), .ZN(p_wishbone_bd_ram_n23785) );
  INV_X1 U32774 ( .A(n62077), .ZN(n28304) );
  INV_X1 U32775 ( .A(n28304), .ZN(p_wishbone_bd_ram_n23784) );
  INV_X1 U32776 ( .A(n62076), .ZN(n28306) );
  INV_X1 U32777 ( .A(n28306), .ZN(p_wishbone_bd_ram_n23783) );
  INV_X1 U32778 ( .A(n62075), .ZN(n28308) );
  INV_X1 U32779 ( .A(n28308), .ZN(p_wishbone_bd_ram_n23782) );
  INV_X1 U32780 ( .A(n62074), .ZN(n28310) );
  INV_X1 U32781 ( .A(n28310), .ZN(p_wishbone_bd_ram_n23781) );
  INV_X1 U32782 ( .A(n62073), .ZN(n28312) );
  INV_X1 U32783 ( .A(n28312), .ZN(p_wishbone_bd_ram_n23780) );
  INV_X1 U32784 ( .A(n62072), .ZN(n28314) );
  INV_X1 U32785 ( .A(n28314), .ZN(p_wishbone_bd_ram_n23779) );
  INV_X1 U32786 ( .A(n62071), .ZN(n28316) );
  INV_X1 U32787 ( .A(n28316), .ZN(p_wishbone_bd_ram_n23778) );
  INV_X1 U32788 ( .A(n62070), .ZN(n28318) );
  INV_X1 U32789 ( .A(n28318), .ZN(p_wishbone_bd_ram_n23777) );
  INV_X1 U32790 ( .A(n62069), .ZN(n28320) );
  INV_X1 U32791 ( .A(n28320), .ZN(p_wishbone_bd_ram_n23776) );
  INV_X1 U32792 ( .A(n62068), .ZN(n28322) );
  INV_X1 U32793 ( .A(n28322), .ZN(p_wishbone_bd_ram_n23775) );
  INV_X1 U32794 ( .A(n62067), .ZN(n28324) );
  INV_X1 U32795 ( .A(n28324), .ZN(p_wishbone_bd_ram_n23774) );
  INV_X1 U32796 ( .A(n62066), .ZN(n28326) );
  INV_X1 U32797 ( .A(n28326), .ZN(p_wishbone_bd_ram_n23773) );
  INV_X1 U32798 ( .A(n62065), .ZN(n28328) );
  INV_X1 U32799 ( .A(n28328), .ZN(p_wishbone_bd_ram_n23772) );
  INV_X1 U32800 ( .A(n62064), .ZN(n28330) );
  INV_X1 U32801 ( .A(n28330), .ZN(p_wishbone_bd_ram_n23771) );
  INV_X1 U32802 ( .A(n62063), .ZN(n28332) );
  INV_X1 U32803 ( .A(n28332), .ZN(p_wishbone_bd_ram_n23770) );
  INV_X1 U32804 ( .A(n62062), .ZN(n28334) );
  INV_X1 U32805 ( .A(n28334), .ZN(p_wishbone_bd_ram_n23769) );
  INV_X1 U32806 ( .A(n62061), .ZN(n28336) );
  INV_X1 U32807 ( .A(n28336), .ZN(p_wishbone_bd_ram_n23768) );
  INV_X1 U32808 ( .A(n62060), .ZN(n28338) );
  INV_X1 U32809 ( .A(n28338), .ZN(p_wishbone_bd_ram_n23767) );
  INV_X1 U32810 ( .A(n62059), .ZN(n28340) );
  INV_X1 U32811 ( .A(n28340), .ZN(p_wishbone_bd_ram_n23766) );
  INV_X1 U32812 ( .A(n62058), .ZN(n28342) );
  INV_X1 U32813 ( .A(n28342), .ZN(p_wishbone_bd_ram_n23765) );
  INV_X1 U32814 ( .A(n62057), .ZN(n28344) );
  INV_X1 U32815 ( .A(n28344), .ZN(p_wishbone_bd_ram_n23764) );
  INV_X1 U32816 ( .A(n62056), .ZN(n28346) );
  INV_X1 U32817 ( .A(n28346), .ZN(p_wishbone_bd_ram_n23763) );
  INV_X1 U32818 ( .A(n62055), .ZN(n28348) );
  INV_X1 U32819 ( .A(n28348), .ZN(p_wishbone_bd_ram_n23762) );
  INV_X1 U32820 ( .A(n62054), .ZN(n28350) );
  INV_X1 U32821 ( .A(n28350), .ZN(p_wishbone_bd_ram_n23761) );
  INV_X1 U32822 ( .A(n62053), .ZN(n28352) );
  INV_X1 U32823 ( .A(n28352), .ZN(p_wishbone_bd_ram_n23760) );
  INV_X1 U32824 ( .A(n62052), .ZN(n28354) );
  INV_X1 U32825 ( .A(n28354), .ZN(p_wishbone_bd_ram_n23759) );
  INV_X1 U32826 ( .A(n62051), .ZN(n28356) );
  INV_X1 U32827 ( .A(n28356), .ZN(p_wishbone_bd_ram_n23758) );
  INV_X1 U32828 ( .A(n62050), .ZN(n28358) );
  INV_X1 U32829 ( .A(n28358), .ZN(p_wishbone_bd_ram_n23757) );
  INV_X1 U32830 ( .A(n62049), .ZN(n28360) );
  INV_X1 U32831 ( .A(n28360), .ZN(p_wishbone_bd_ram_n23756) );
  INV_X1 U32832 ( .A(n62048), .ZN(n28362) );
  INV_X1 U32833 ( .A(n28362), .ZN(p_wishbone_bd_ram_n23755) );
  INV_X1 U32834 ( .A(n62047), .ZN(n28364) );
  INV_X1 U32835 ( .A(n28364), .ZN(p_wishbone_bd_ram_n23754) );
  INV_X1 U32836 ( .A(n62046), .ZN(n28366) );
  INV_X1 U32837 ( .A(n28366), .ZN(p_wishbone_bd_ram_n23753) );
  INV_X1 U32838 ( .A(n62045), .ZN(n28368) );
  INV_X1 U32839 ( .A(n28368), .ZN(p_wishbone_bd_ram_n23752) );
  INV_X1 U32840 ( .A(n62044), .ZN(n28370) );
  INV_X1 U32841 ( .A(n28370), .ZN(p_wishbone_bd_ram_n23751) );
  INV_X1 U32842 ( .A(n62043), .ZN(n28372) );
  INV_X1 U32843 ( .A(n28372), .ZN(p_wishbone_bd_ram_n23750) );
  INV_X1 U32844 ( .A(n62042), .ZN(n28374) );
  INV_X1 U32845 ( .A(n28374), .ZN(p_wishbone_bd_ram_n23749) );
  INV_X1 U32846 ( .A(n62041), .ZN(n28376) );
  INV_X1 U32847 ( .A(n28376), .ZN(p_wishbone_bd_ram_n23748) );
  INV_X1 U32848 ( .A(n62040), .ZN(n28378) );
  INV_X1 U32849 ( .A(n28378), .ZN(p_wishbone_bd_ram_n23747) );
  INV_X1 U32850 ( .A(n62039), .ZN(n28380) );
  INV_X1 U32851 ( .A(n28380), .ZN(p_wishbone_bd_ram_n23746) );
  INV_X1 U32852 ( .A(n62038), .ZN(n28382) );
  INV_X1 U32853 ( .A(n28382), .ZN(p_wishbone_bd_ram_n23745) );
  INV_X1 U32854 ( .A(n62037), .ZN(n28384) );
  INV_X1 U32855 ( .A(n28384), .ZN(p_wishbone_bd_ram_n23744) );
  INV_X1 U32856 ( .A(n62036), .ZN(n28386) );
  INV_X1 U32857 ( .A(n28386), .ZN(p_wishbone_bd_ram_n23743) );
  INV_X1 U32858 ( .A(n62035), .ZN(n28388) );
  INV_X1 U32859 ( .A(n28388), .ZN(p_wishbone_bd_ram_n23742) );
  INV_X1 U32860 ( .A(n62034), .ZN(n28390) );
  INV_X1 U32861 ( .A(n28390), .ZN(p_wishbone_bd_ram_n23741) );
  INV_X1 U32862 ( .A(n62033), .ZN(n28392) );
  INV_X1 U32863 ( .A(n28392), .ZN(p_wishbone_bd_ram_n23740) );
  INV_X1 U32864 ( .A(n62032), .ZN(n28394) );
  INV_X1 U32865 ( .A(n28394), .ZN(p_wishbone_bd_ram_n23739) );
  INV_X1 U32866 ( .A(n62031), .ZN(n28396) );
  INV_X1 U32867 ( .A(n28396), .ZN(p_wishbone_bd_ram_n23738) );
  INV_X1 U32868 ( .A(n62030), .ZN(n28398) );
  INV_X1 U32869 ( .A(n28398), .ZN(p_wishbone_bd_ram_n23737) );
  INV_X1 U32870 ( .A(n62029), .ZN(n28400) );
  INV_X1 U32871 ( .A(n28400), .ZN(p_wishbone_bd_ram_n23736) );
  INV_X1 U32872 ( .A(n62028), .ZN(n28402) );
  INV_X1 U32873 ( .A(n28402), .ZN(p_wishbone_bd_ram_n23735) );
  INV_X1 U32874 ( .A(n62027), .ZN(n28404) );
  INV_X1 U32875 ( .A(n28404), .ZN(p_wishbone_bd_ram_n23734) );
  INV_X1 U32876 ( .A(n62026), .ZN(n28406) );
  INV_X1 U32877 ( .A(n28406), .ZN(p_wishbone_bd_ram_n23733) );
  INV_X1 U32878 ( .A(n62025), .ZN(n28408) );
  INV_X1 U32879 ( .A(n28408), .ZN(p_wishbone_bd_ram_n23732) );
  INV_X1 U32880 ( .A(n62024), .ZN(n28410) );
  INV_X1 U32881 ( .A(n28410), .ZN(p_wishbone_bd_ram_n23731) );
  INV_X1 U32882 ( .A(n62023), .ZN(n28412) );
  INV_X1 U32883 ( .A(n28412), .ZN(p_wishbone_bd_ram_n23730) );
  INV_X1 U32884 ( .A(n62022), .ZN(n28414) );
  INV_X1 U32885 ( .A(n28414), .ZN(p_wishbone_bd_ram_n23729) );
  INV_X1 U32886 ( .A(n62021), .ZN(n28416) );
  INV_X1 U32887 ( .A(n28416), .ZN(p_wishbone_bd_ram_n23728) );
  INV_X1 U32888 ( .A(n62020), .ZN(n28418) );
  INV_X1 U32889 ( .A(n28418), .ZN(p_wishbone_bd_ram_n23727) );
  INV_X1 U32890 ( .A(n62019), .ZN(n28420) );
  INV_X1 U32891 ( .A(n28420), .ZN(p_wishbone_bd_ram_n23726) );
  INV_X1 U32892 ( .A(n62018), .ZN(n28422) );
  INV_X1 U32893 ( .A(n28422), .ZN(p_wishbone_bd_ram_n23725) );
  INV_X1 U32894 ( .A(n62017), .ZN(n28424) );
  INV_X1 U32895 ( .A(n28424), .ZN(p_wishbone_bd_ram_n23724) );
  INV_X1 U32896 ( .A(n62016), .ZN(n28426) );
  INV_X1 U32897 ( .A(n28426), .ZN(p_wishbone_bd_ram_n23723) );
  INV_X1 U32898 ( .A(n62015), .ZN(n28428) );
  INV_X1 U32899 ( .A(n28428), .ZN(p_wishbone_bd_ram_n23722) );
  INV_X1 U32900 ( .A(n62014), .ZN(n28430) );
  INV_X1 U32901 ( .A(n28430), .ZN(p_wishbone_bd_ram_n23721) );
  INV_X1 U32902 ( .A(n62013), .ZN(n28432) );
  INV_X1 U32903 ( .A(n28432), .ZN(p_wishbone_bd_ram_n23720) );
  INV_X1 U32904 ( .A(n62012), .ZN(n28434) );
  INV_X1 U32905 ( .A(n28434), .ZN(p_wishbone_bd_ram_n23719) );
  INV_X1 U32906 ( .A(n62011), .ZN(n28436) );
  INV_X1 U32907 ( .A(n28436), .ZN(p_wishbone_bd_ram_n23718) );
  INV_X1 U32908 ( .A(n62010), .ZN(n28438) );
  INV_X1 U32909 ( .A(n28438), .ZN(p_wishbone_bd_ram_n23717) );
  INV_X1 U32910 ( .A(n62009), .ZN(n28440) );
  INV_X1 U32911 ( .A(n28440), .ZN(p_wishbone_bd_ram_n23716) );
  INV_X1 U32912 ( .A(n62008), .ZN(n28442) );
  INV_X1 U32913 ( .A(n28442), .ZN(p_wishbone_bd_ram_n23715) );
  INV_X1 U32914 ( .A(n62007), .ZN(n28444) );
  INV_X1 U32915 ( .A(n28444), .ZN(p_wishbone_bd_ram_n23714) );
  INV_X1 U32916 ( .A(n62006), .ZN(n28446) );
  INV_X1 U32917 ( .A(n28446), .ZN(p_wishbone_bd_ram_n23713) );
  INV_X1 U32918 ( .A(n62005), .ZN(n28448) );
  INV_X1 U32919 ( .A(n28448), .ZN(p_wishbone_bd_ram_n23712) );
  INV_X1 U32920 ( .A(n62004), .ZN(n28450) );
  INV_X1 U32921 ( .A(n28450), .ZN(p_wishbone_bd_ram_n23711) );
  INV_X1 U32922 ( .A(n62003), .ZN(n28452) );
  INV_X1 U32923 ( .A(n28452), .ZN(p_wishbone_bd_ram_n23710) );
  INV_X1 U32924 ( .A(n62002), .ZN(n28454) );
  INV_X1 U32925 ( .A(n28454), .ZN(p_wishbone_bd_ram_n23709) );
  INV_X1 U32926 ( .A(n62001), .ZN(n28456) );
  INV_X1 U32927 ( .A(n28456), .ZN(p_wishbone_bd_ram_n23708) );
  INV_X1 U32928 ( .A(n62000), .ZN(n28458) );
  INV_X1 U32929 ( .A(n28458), .ZN(p_wishbone_bd_ram_n23707) );
  INV_X1 U32930 ( .A(n61999), .ZN(n28460) );
  INV_X1 U32931 ( .A(n28460), .ZN(p_wishbone_bd_ram_n23706) );
  INV_X1 U32932 ( .A(n61998), .ZN(n28462) );
  INV_X1 U32933 ( .A(n28462), .ZN(p_wishbone_bd_ram_n23705) );
  INV_X1 U32934 ( .A(n61997), .ZN(n28464) );
  INV_X1 U32935 ( .A(n28464), .ZN(p_wishbone_bd_ram_n23704) );
  INV_X1 U32936 ( .A(n61996), .ZN(n28466) );
  INV_X1 U32937 ( .A(n28466), .ZN(p_wishbone_bd_ram_n23703) );
  INV_X1 U32938 ( .A(n61995), .ZN(n28468) );
  INV_X1 U32939 ( .A(n28468), .ZN(p_wishbone_bd_ram_n23702) );
  INV_X1 U32940 ( .A(n61994), .ZN(n28470) );
  INV_X1 U32941 ( .A(n28470), .ZN(p_wishbone_bd_ram_n23701) );
  INV_X1 U32942 ( .A(n61993), .ZN(n28472) );
  INV_X1 U32943 ( .A(n28472), .ZN(p_wishbone_bd_ram_n23700) );
  INV_X1 U32944 ( .A(n61992), .ZN(n28474) );
  INV_X1 U32945 ( .A(n28474), .ZN(p_wishbone_bd_ram_n23699) );
  INV_X1 U32946 ( .A(n61991), .ZN(n28476) );
  INV_X1 U32947 ( .A(n28476), .ZN(p_wishbone_bd_ram_n23698) );
  INV_X1 U32948 ( .A(n61990), .ZN(n28478) );
  INV_X1 U32949 ( .A(n28478), .ZN(p_wishbone_bd_ram_n23697) );
  INV_X1 U32950 ( .A(n61989), .ZN(n28480) );
  INV_X1 U32951 ( .A(n28480), .ZN(p_wishbone_bd_ram_n23696) );
  INV_X1 U32952 ( .A(n61988), .ZN(n28482) );
  INV_X1 U32953 ( .A(n28482), .ZN(p_wishbone_bd_ram_n23695) );
  INV_X1 U32954 ( .A(n61987), .ZN(n28484) );
  INV_X1 U32955 ( .A(n28484), .ZN(p_wishbone_bd_ram_n23694) );
  INV_X1 U32956 ( .A(n61986), .ZN(n28486) );
  INV_X1 U32957 ( .A(n28486), .ZN(p_wishbone_bd_ram_n23693) );
  INV_X1 U32958 ( .A(n61985), .ZN(n28488) );
  INV_X1 U32959 ( .A(n28488), .ZN(p_wishbone_bd_ram_n23692) );
  INV_X1 U32960 ( .A(n61984), .ZN(n28490) );
  INV_X1 U32961 ( .A(n28490), .ZN(p_wishbone_bd_ram_n23691) );
  INV_X1 U32962 ( .A(n61983), .ZN(n28492) );
  INV_X1 U32963 ( .A(n28492), .ZN(p_wishbone_bd_ram_n23690) );
  INV_X1 U32964 ( .A(n61982), .ZN(n28494) );
  INV_X1 U32965 ( .A(n28494), .ZN(p_wishbone_bd_ram_n23689) );
  INV_X1 U32966 ( .A(n61981), .ZN(n28496) );
  INV_X1 U32967 ( .A(n28496), .ZN(p_wishbone_bd_ram_n23688) );
  INV_X1 U32968 ( .A(n61980), .ZN(n28498) );
  INV_X1 U32969 ( .A(n28498), .ZN(p_wishbone_bd_ram_n23687) );
  INV_X1 U32970 ( .A(n61979), .ZN(n28500) );
  INV_X1 U32971 ( .A(n28500), .ZN(p_wishbone_bd_ram_n23686) );
  INV_X1 U32972 ( .A(n61978), .ZN(n28502) );
  INV_X1 U32973 ( .A(n28502), .ZN(p_wishbone_bd_ram_n23685) );
  INV_X1 U32974 ( .A(n61977), .ZN(n28504) );
  INV_X1 U32975 ( .A(n28504), .ZN(p_wishbone_bd_ram_n23684) );
  INV_X1 U32976 ( .A(n61976), .ZN(n28506) );
  INV_X1 U32977 ( .A(n28506), .ZN(p_wishbone_bd_ram_n23683) );
  INV_X1 U32978 ( .A(n61975), .ZN(n28508) );
  INV_X1 U32979 ( .A(n28508), .ZN(p_wishbone_bd_ram_n23682) );
  INV_X1 U32980 ( .A(n61974), .ZN(n28510) );
  INV_X1 U32981 ( .A(n28510), .ZN(p_wishbone_bd_ram_n23681) );
  INV_X1 U32982 ( .A(n61973), .ZN(n28512) );
  INV_X1 U32983 ( .A(n28512), .ZN(p_wishbone_bd_ram_n23680) );
  INV_X1 U32984 ( .A(n61972), .ZN(n28514) );
  INV_X1 U32985 ( .A(n28514), .ZN(p_wishbone_bd_ram_n23679) );
  INV_X1 U32986 ( .A(n61971), .ZN(n28516) );
  INV_X1 U32987 ( .A(n28516), .ZN(p_wishbone_bd_ram_n23678) );
  INV_X1 U32988 ( .A(n61970), .ZN(n28518) );
  INV_X1 U32989 ( .A(n28518), .ZN(p_wishbone_bd_ram_n23677) );
  INV_X1 U32990 ( .A(n61969), .ZN(n28520) );
  INV_X1 U32991 ( .A(n28520), .ZN(p_wishbone_bd_ram_n23676) );
  INV_X1 U32992 ( .A(n61968), .ZN(n28522) );
  INV_X1 U32993 ( .A(n28522), .ZN(p_wishbone_bd_ram_n23675) );
  INV_X1 U32994 ( .A(n61967), .ZN(n28524) );
  INV_X1 U32995 ( .A(n28524), .ZN(p_wishbone_bd_ram_n23674) );
  INV_X1 U32996 ( .A(n61966), .ZN(n28526) );
  INV_X1 U32997 ( .A(n28526), .ZN(p_wishbone_bd_ram_n23673) );
  INV_X1 U32998 ( .A(n61965), .ZN(n28528) );
  INV_X1 U32999 ( .A(n28528), .ZN(p_wishbone_bd_ram_n23672) );
  INV_X1 U33000 ( .A(n61964), .ZN(n28530) );
  INV_X1 U33001 ( .A(n28530), .ZN(p_wishbone_bd_ram_n23671) );
  INV_X1 U33002 ( .A(n61963), .ZN(n28532) );
  INV_X1 U33003 ( .A(n28532), .ZN(p_wishbone_bd_ram_n23670) );
  INV_X1 U33004 ( .A(n61962), .ZN(n28534) );
  INV_X1 U33005 ( .A(n28534), .ZN(p_wishbone_bd_ram_n23669) );
  INV_X1 U33006 ( .A(n61961), .ZN(n28536) );
  INV_X1 U33007 ( .A(n28536), .ZN(p_wishbone_bd_ram_n23668) );
  INV_X1 U33008 ( .A(n61960), .ZN(n28538) );
  INV_X1 U33009 ( .A(n28538), .ZN(p_wishbone_bd_ram_n23667) );
  INV_X1 U33010 ( .A(n61959), .ZN(n28540) );
  INV_X1 U33011 ( .A(n28540), .ZN(p_wishbone_bd_ram_n23666) );
  INV_X1 U33012 ( .A(n61958), .ZN(n28542) );
  INV_X1 U33013 ( .A(n28542), .ZN(p_wishbone_bd_ram_n23665) );
  INV_X1 U33014 ( .A(n61957), .ZN(n28544) );
  INV_X1 U33015 ( .A(n28544), .ZN(p_wishbone_bd_ram_n23664) );
  INV_X1 U33016 ( .A(n61956), .ZN(n28546) );
  INV_X1 U33017 ( .A(n28546), .ZN(p_wishbone_bd_ram_n23663) );
  INV_X1 U33018 ( .A(n61955), .ZN(n28548) );
  INV_X1 U33019 ( .A(n28548), .ZN(p_wishbone_bd_ram_n23662) );
  INV_X1 U33020 ( .A(n61954), .ZN(n28550) );
  INV_X1 U33021 ( .A(n28550), .ZN(p_wishbone_bd_ram_n23661) );
  INV_X1 U33022 ( .A(n61953), .ZN(n28552) );
  INV_X1 U33023 ( .A(n28552), .ZN(p_wishbone_bd_ram_n23660) );
  INV_X1 U33024 ( .A(n61952), .ZN(n28554) );
  INV_X1 U33025 ( .A(n28554), .ZN(p_wishbone_bd_ram_n23659) );
  INV_X1 U33026 ( .A(n61951), .ZN(n28556) );
  INV_X1 U33027 ( .A(n28556), .ZN(p_wishbone_bd_ram_n23658) );
  INV_X1 U33028 ( .A(n61950), .ZN(n28558) );
  INV_X1 U33029 ( .A(n28558), .ZN(p_wishbone_bd_ram_n23657) );
  INV_X1 U33030 ( .A(n61949), .ZN(n28560) );
  INV_X1 U33031 ( .A(n28560), .ZN(p_wishbone_bd_ram_n23656) );
  INV_X1 U33032 ( .A(n61948), .ZN(n28562) );
  INV_X1 U33033 ( .A(n28562), .ZN(p_wishbone_bd_ram_n23655) );
  INV_X1 U33034 ( .A(n61947), .ZN(n28564) );
  INV_X1 U33035 ( .A(n28564), .ZN(p_wishbone_bd_ram_n23654) );
  INV_X1 U33036 ( .A(n61946), .ZN(n28566) );
  INV_X1 U33037 ( .A(n28566), .ZN(p_wishbone_bd_ram_n23653) );
  INV_X1 U33038 ( .A(n61945), .ZN(n28568) );
  INV_X1 U33039 ( .A(n28568), .ZN(p_wishbone_bd_ram_n23652) );
  INV_X1 U33040 ( .A(n61944), .ZN(n28570) );
  INV_X1 U33041 ( .A(n28570), .ZN(p_wishbone_bd_ram_n23651) );
  INV_X1 U33042 ( .A(n61943), .ZN(n28572) );
  INV_X1 U33043 ( .A(n28572), .ZN(p_wishbone_bd_ram_n23650) );
  INV_X1 U33044 ( .A(n61942), .ZN(n28574) );
  INV_X1 U33045 ( .A(n28574), .ZN(p_wishbone_bd_ram_n23649) );
  INV_X1 U33046 ( .A(n61941), .ZN(n28576) );
  INV_X1 U33047 ( .A(n28576), .ZN(p_wishbone_bd_ram_n23648) );
  INV_X1 U33048 ( .A(n61940), .ZN(n28578) );
  INV_X1 U33049 ( .A(n28578), .ZN(p_wishbone_bd_ram_n23647) );
  INV_X1 U33050 ( .A(n61939), .ZN(n28580) );
  INV_X1 U33051 ( .A(n28580), .ZN(p_wishbone_bd_ram_n23646) );
  INV_X1 U33052 ( .A(n61938), .ZN(n28582) );
  INV_X1 U33053 ( .A(n28582), .ZN(p_wishbone_bd_ram_n23645) );
  INV_X1 U33054 ( .A(n61937), .ZN(n28584) );
  INV_X1 U33055 ( .A(n28584), .ZN(p_wishbone_bd_ram_n23644) );
  INV_X1 U33056 ( .A(n61936), .ZN(n28586) );
  INV_X1 U33057 ( .A(n28586), .ZN(p_wishbone_bd_ram_n23643) );
  INV_X1 U33058 ( .A(n61935), .ZN(n28588) );
  INV_X1 U33059 ( .A(n28588), .ZN(p_wishbone_bd_ram_n23642) );
  INV_X1 U33060 ( .A(n61934), .ZN(n28590) );
  INV_X1 U33061 ( .A(n28590), .ZN(p_wishbone_bd_ram_n23641) );
  INV_X1 U33062 ( .A(n61933), .ZN(n28592) );
  INV_X1 U33063 ( .A(n28592), .ZN(p_wishbone_bd_ram_n23640) );
  INV_X1 U33064 ( .A(n61932), .ZN(n28594) );
  INV_X1 U33065 ( .A(n28594), .ZN(p_wishbone_bd_ram_n23639) );
  INV_X1 U33066 ( .A(n61931), .ZN(n28596) );
  INV_X1 U33067 ( .A(n28596), .ZN(p_wishbone_bd_ram_n23638) );
  INV_X1 U33068 ( .A(n61930), .ZN(n28598) );
  INV_X1 U33069 ( .A(n28598), .ZN(p_wishbone_bd_ram_n23637) );
  INV_X1 U33070 ( .A(n61929), .ZN(n28600) );
  INV_X1 U33071 ( .A(n28600), .ZN(p_wishbone_bd_ram_n23636) );
  INV_X1 U33072 ( .A(n61928), .ZN(n28602) );
  INV_X1 U33073 ( .A(n28602), .ZN(p_wishbone_bd_ram_n23635) );
  INV_X1 U33074 ( .A(n61927), .ZN(n28604) );
  INV_X1 U33075 ( .A(n28604), .ZN(p_wishbone_bd_ram_n23634) );
  INV_X1 U33076 ( .A(n61926), .ZN(n28606) );
  INV_X1 U33077 ( .A(n28606), .ZN(p_wishbone_bd_ram_n23633) );
  INV_X1 U33078 ( .A(n61925), .ZN(n28608) );
  INV_X1 U33079 ( .A(n28608), .ZN(p_wishbone_bd_ram_n23632) );
  INV_X1 U33080 ( .A(n61924), .ZN(n28610) );
  INV_X1 U33081 ( .A(n28610), .ZN(p_wishbone_bd_ram_n23631) );
  INV_X1 U33082 ( .A(n61923), .ZN(n28612) );
  INV_X1 U33083 ( .A(n28612), .ZN(p_wishbone_bd_ram_n23630) );
  INV_X1 U33084 ( .A(n61922), .ZN(n28614) );
  INV_X1 U33085 ( .A(n28614), .ZN(p_wishbone_bd_ram_n23629) );
  INV_X1 U33086 ( .A(n61921), .ZN(n28616) );
  INV_X1 U33087 ( .A(n28616), .ZN(p_wishbone_bd_ram_n23628) );
  INV_X1 U33088 ( .A(n61920), .ZN(n28618) );
  INV_X1 U33089 ( .A(n28618), .ZN(p_wishbone_bd_ram_n23627) );
  INV_X1 U33090 ( .A(n61919), .ZN(n28620) );
  INV_X1 U33091 ( .A(n28620), .ZN(p_wishbone_bd_ram_n23626) );
  INV_X1 U33092 ( .A(n61918), .ZN(n28622) );
  INV_X1 U33093 ( .A(n28622), .ZN(p_wishbone_bd_ram_n23625) );
  INV_X1 U33094 ( .A(n61917), .ZN(n28624) );
  INV_X1 U33095 ( .A(n28624), .ZN(p_wishbone_bd_ram_n23624) );
  INV_X1 U33096 ( .A(n61916), .ZN(n28626) );
  INV_X1 U33097 ( .A(n28626), .ZN(p_wishbone_bd_ram_n23623) );
  INV_X1 U33098 ( .A(n61915), .ZN(n28628) );
  INV_X1 U33099 ( .A(n28628), .ZN(p_wishbone_bd_ram_n23622) );
  INV_X1 U33100 ( .A(n61914), .ZN(n28630) );
  INV_X1 U33101 ( .A(n28630), .ZN(p_wishbone_bd_ram_n23621) );
  INV_X1 U33102 ( .A(n61913), .ZN(n28632) );
  INV_X1 U33103 ( .A(n28632), .ZN(p_wishbone_bd_ram_n23620) );
  INV_X1 U33104 ( .A(n61912), .ZN(n28634) );
  INV_X1 U33105 ( .A(n28634), .ZN(p_wishbone_bd_ram_n23619) );
  INV_X1 U33106 ( .A(n61911), .ZN(n28636) );
  INV_X1 U33107 ( .A(n28636), .ZN(p_wishbone_bd_ram_n23618) );
  INV_X1 U33108 ( .A(n61910), .ZN(n28638) );
  INV_X1 U33109 ( .A(n28638), .ZN(p_wishbone_bd_ram_n23617) );
  INV_X1 U33110 ( .A(n61909), .ZN(n28640) );
  INV_X1 U33111 ( .A(n28640), .ZN(p_wishbone_bd_ram_n23616) );
  INV_X1 U33112 ( .A(n61908), .ZN(n28642) );
  INV_X1 U33113 ( .A(n28642), .ZN(p_wishbone_bd_ram_n23615) );
  INV_X1 U33114 ( .A(n61907), .ZN(n28644) );
  INV_X1 U33115 ( .A(n28644), .ZN(p_wishbone_bd_ram_n23614) );
  INV_X1 U33116 ( .A(n61906), .ZN(n28646) );
  INV_X1 U33117 ( .A(n28646), .ZN(p_wishbone_bd_ram_n23613) );
  INV_X1 U33118 ( .A(n61905), .ZN(n28648) );
  INV_X1 U33119 ( .A(n28648), .ZN(p_wishbone_bd_ram_n23612) );
  INV_X1 U33120 ( .A(n61904), .ZN(n28650) );
  INV_X1 U33121 ( .A(n28650), .ZN(p_wishbone_bd_ram_n23611) );
  INV_X1 U33122 ( .A(n61903), .ZN(n28652) );
  INV_X1 U33123 ( .A(n28652), .ZN(p_wishbone_bd_ram_n23610) );
  INV_X1 U33124 ( .A(n61902), .ZN(n28654) );
  INV_X1 U33125 ( .A(n28654), .ZN(p_wishbone_bd_ram_n23609) );
  INV_X1 U33126 ( .A(n61901), .ZN(n28656) );
  INV_X1 U33127 ( .A(n28656), .ZN(p_wishbone_bd_ram_n23608) );
  INV_X1 U33128 ( .A(n61900), .ZN(n28658) );
  INV_X1 U33129 ( .A(n28658), .ZN(p_wishbone_bd_ram_n23607) );
  INV_X1 U33130 ( .A(n61899), .ZN(n28660) );
  INV_X1 U33131 ( .A(n28660), .ZN(p_wishbone_bd_ram_n23606) );
  INV_X1 U33132 ( .A(n61898), .ZN(n28662) );
  INV_X1 U33133 ( .A(n28662), .ZN(p_wishbone_bd_ram_n23605) );
  INV_X1 U33134 ( .A(n61897), .ZN(n28664) );
  INV_X1 U33135 ( .A(n28664), .ZN(p_wishbone_bd_ram_n23604) );
  INV_X1 U33136 ( .A(n61896), .ZN(n28666) );
  INV_X1 U33137 ( .A(n28666), .ZN(p_wishbone_bd_ram_n23603) );
  INV_X1 U33138 ( .A(n61895), .ZN(n28668) );
  INV_X1 U33139 ( .A(n28668), .ZN(p_wishbone_bd_ram_n23602) );
  INV_X1 U33140 ( .A(n61894), .ZN(n28670) );
  INV_X1 U33141 ( .A(n28670), .ZN(p_wishbone_bd_ram_n23601) );
  INV_X1 U33142 ( .A(n61893), .ZN(n28672) );
  INV_X1 U33143 ( .A(n28672), .ZN(p_wishbone_bd_ram_n23600) );
  INV_X1 U33144 ( .A(n61892), .ZN(n28674) );
  INV_X1 U33145 ( .A(n28674), .ZN(p_wishbone_bd_ram_n23599) );
  INV_X1 U33146 ( .A(n61891), .ZN(n28676) );
  INV_X1 U33147 ( .A(n28676), .ZN(p_wishbone_bd_ram_n23598) );
  INV_X1 U33148 ( .A(n61890), .ZN(n28678) );
  INV_X1 U33149 ( .A(n28678), .ZN(p_wishbone_bd_ram_n23597) );
  INV_X1 U33150 ( .A(n61889), .ZN(n28680) );
  INV_X1 U33151 ( .A(n28680), .ZN(p_wishbone_bd_ram_n23596) );
  INV_X1 U33152 ( .A(n61888), .ZN(n28682) );
  INV_X1 U33153 ( .A(n28682), .ZN(p_wishbone_bd_ram_n23595) );
  INV_X1 U33154 ( .A(n61887), .ZN(n28684) );
  INV_X1 U33155 ( .A(n28684), .ZN(p_wishbone_bd_ram_n23594) );
  INV_X1 U33156 ( .A(n61886), .ZN(n28686) );
  INV_X1 U33157 ( .A(n28686), .ZN(p_wishbone_bd_ram_n23593) );
  INV_X1 U33158 ( .A(n61885), .ZN(n28688) );
  INV_X1 U33159 ( .A(n28688), .ZN(p_wishbone_bd_ram_n23592) );
  INV_X1 U33160 ( .A(n61884), .ZN(n28690) );
  INV_X1 U33161 ( .A(n28690), .ZN(p_wishbone_bd_ram_n23591) );
  INV_X1 U33162 ( .A(n61883), .ZN(n28692) );
  INV_X1 U33163 ( .A(n28692), .ZN(p_wishbone_bd_ram_n23590) );
  INV_X1 U33164 ( .A(n61882), .ZN(n28694) );
  INV_X1 U33165 ( .A(n28694), .ZN(p_wishbone_bd_ram_n23589) );
  INV_X1 U33166 ( .A(n61881), .ZN(n28696) );
  INV_X1 U33167 ( .A(n28696), .ZN(p_wishbone_bd_ram_n23588) );
  INV_X1 U33168 ( .A(n61880), .ZN(n28698) );
  INV_X1 U33169 ( .A(n28698), .ZN(p_wishbone_bd_ram_n23587) );
  INV_X1 U33170 ( .A(n61879), .ZN(n28700) );
  INV_X1 U33171 ( .A(n28700), .ZN(p_wishbone_bd_ram_n23586) );
  INV_X1 U33172 ( .A(n61878), .ZN(n28702) );
  INV_X1 U33173 ( .A(n28702), .ZN(p_wishbone_bd_ram_n23585) );
  INV_X1 U33174 ( .A(n61877), .ZN(n28704) );
  INV_X1 U33175 ( .A(n28704), .ZN(p_wishbone_bd_ram_n23584) );
  INV_X1 U33176 ( .A(n61876), .ZN(n28706) );
  INV_X1 U33177 ( .A(n28706), .ZN(p_wishbone_bd_ram_n23583) );
  INV_X1 U33178 ( .A(n61875), .ZN(n28708) );
  INV_X1 U33179 ( .A(n28708), .ZN(p_wishbone_bd_ram_n23582) );
  INV_X1 U33180 ( .A(n61874), .ZN(n28710) );
  INV_X1 U33181 ( .A(n28710), .ZN(p_wishbone_bd_ram_n23581) );
  INV_X1 U33182 ( .A(n61873), .ZN(n28712) );
  INV_X1 U33183 ( .A(n28712), .ZN(p_wishbone_bd_ram_n23580) );
  INV_X1 U33184 ( .A(n61872), .ZN(n28714) );
  INV_X1 U33185 ( .A(n28714), .ZN(p_wishbone_bd_ram_n23579) );
  INV_X1 U33186 ( .A(n61871), .ZN(n28716) );
  INV_X1 U33187 ( .A(n28716), .ZN(p_wishbone_bd_ram_n23578) );
  INV_X1 U33188 ( .A(n61870), .ZN(n28718) );
  INV_X1 U33189 ( .A(n28718), .ZN(p_wishbone_bd_ram_n23577) );
  INV_X1 U33190 ( .A(n61869), .ZN(n28720) );
  INV_X1 U33191 ( .A(n28720), .ZN(p_wishbone_bd_ram_n23576) );
  INV_X1 U33192 ( .A(n61868), .ZN(n28722) );
  INV_X1 U33193 ( .A(n28722), .ZN(p_wishbone_bd_ram_n23575) );
  INV_X1 U33194 ( .A(n61867), .ZN(n28724) );
  INV_X1 U33195 ( .A(n28724), .ZN(p_wishbone_bd_ram_n23574) );
  INV_X1 U33196 ( .A(n61866), .ZN(n28726) );
  INV_X1 U33197 ( .A(n28726), .ZN(p_wishbone_bd_ram_n23573) );
  INV_X1 U33198 ( .A(n61865), .ZN(n28728) );
  INV_X1 U33199 ( .A(n28728), .ZN(p_wishbone_bd_ram_n23572) );
  INV_X1 U33200 ( .A(n61864), .ZN(n28730) );
  INV_X1 U33201 ( .A(n28730), .ZN(p_wishbone_bd_ram_n23571) );
  INV_X1 U33202 ( .A(n61863), .ZN(n28732) );
  INV_X1 U33203 ( .A(n28732), .ZN(p_wishbone_bd_ram_n23570) );
  INV_X1 U33204 ( .A(n61862), .ZN(n28734) );
  INV_X1 U33205 ( .A(n28734), .ZN(p_wishbone_bd_ram_n23569) );
  INV_X1 U33206 ( .A(n61861), .ZN(n28736) );
  INV_X1 U33207 ( .A(n28736), .ZN(p_wishbone_bd_ram_n23568) );
  INV_X1 U33208 ( .A(n61860), .ZN(n28738) );
  INV_X1 U33209 ( .A(n28738), .ZN(p_wishbone_bd_ram_n23567) );
  INV_X1 U33210 ( .A(n61859), .ZN(n28740) );
  INV_X1 U33211 ( .A(n28740), .ZN(p_wishbone_bd_ram_n23566) );
  INV_X1 U33212 ( .A(n61858), .ZN(n28742) );
  INV_X1 U33213 ( .A(n28742), .ZN(p_wishbone_bd_ram_n23565) );
  INV_X1 U33214 ( .A(n61857), .ZN(n28744) );
  INV_X1 U33215 ( .A(n28744), .ZN(p_wishbone_bd_ram_n23564) );
  INV_X1 U33216 ( .A(n61856), .ZN(n28746) );
  INV_X1 U33217 ( .A(n28746), .ZN(p_wishbone_bd_ram_n23563) );
  INV_X1 U33218 ( .A(n61855), .ZN(n28748) );
  INV_X1 U33219 ( .A(n28748), .ZN(p_wishbone_bd_ram_n23562) );
  INV_X1 U33220 ( .A(n61854), .ZN(n28750) );
  INV_X1 U33221 ( .A(n28750), .ZN(p_wishbone_bd_ram_n23561) );
  INV_X1 U33222 ( .A(n61853), .ZN(n28752) );
  INV_X1 U33223 ( .A(n28752), .ZN(p_wishbone_bd_ram_n23560) );
  INV_X1 U33224 ( .A(n61852), .ZN(n28754) );
  INV_X1 U33225 ( .A(n28754), .ZN(p_wishbone_bd_ram_n23559) );
  INV_X1 U33226 ( .A(n61851), .ZN(n28756) );
  INV_X1 U33227 ( .A(n28756), .ZN(p_wishbone_bd_ram_n23558) );
  INV_X1 U33228 ( .A(n61850), .ZN(n28758) );
  INV_X1 U33229 ( .A(n28758), .ZN(p_wishbone_bd_ram_n23557) );
  INV_X1 U33230 ( .A(n61849), .ZN(n28760) );
  INV_X1 U33231 ( .A(n28760), .ZN(p_wishbone_bd_ram_n23556) );
  INV_X1 U33232 ( .A(n61848), .ZN(n28762) );
  INV_X1 U33233 ( .A(n28762), .ZN(p_wishbone_bd_ram_n23555) );
  INV_X1 U33234 ( .A(n61847), .ZN(n28764) );
  INV_X1 U33235 ( .A(n28764), .ZN(p_wishbone_bd_ram_n23554) );
  INV_X1 U33236 ( .A(n61846), .ZN(n28766) );
  INV_X1 U33237 ( .A(n28766), .ZN(p_wishbone_bd_ram_n23553) );
  INV_X1 U33238 ( .A(n61845), .ZN(n28768) );
  INV_X1 U33239 ( .A(n28768), .ZN(p_wishbone_bd_ram_n23552) );
  INV_X1 U33240 ( .A(n61844), .ZN(n28770) );
  INV_X1 U33241 ( .A(n28770), .ZN(p_wishbone_bd_ram_n23551) );
  INV_X1 U33242 ( .A(n61843), .ZN(n28772) );
  INV_X1 U33243 ( .A(n28772), .ZN(p_wishbone_bd_ram_n23550) );
  INV_X1 U33244 ( .A(n61842), .ZN(n28774) );
  INV_X1 U33245 ( .A(n28774), .ZN(p_wishbone_bd_ram_n23549) );
  INV_X1 U33246 ( .A(n61841), .ZN(n28776) );
  INV_X1 U33247 ( .A(n28776), .ZN(p_wishbone_bd_ram_n23548) );
  INV_X1 U33248 ( .A(n61840), .ZN(n28778) );
  INV_X1 U33249 ( .A(n28778), .ZN(p_wishbone_bd_ram_n23547) );
  INV_X1 U33250 ( .A(n61839), .ZN(n28780) );
  INV_X1 U33251 ( .A(n28780), .ZN(p_wishbone_bd_ram_n23546) );
  INV_X1 U33252 ( .A(n61838), .ZN(n28782) );
  INV_X1 U33253 ( .A(n28782), .ZN(p_wishbone_bd_ram_n23545) );
  INV_X1 U33254 ( .A(n61837), .ZN(n28784) );
  INV_X1 U33255 ( .A(n28784), .ZN(p_wishbone_bd_ram_n23544) );
  INV_X1 U33256 ( .A(n61836), .ZN(n28786) );
  INV_X1 U33257 ( .A(n28786), .ZN(p_wishbone_bd_ram_n23543) );
  INV_X1 U33258 ( .A(n61835), .ZN(n28788) );
  INV_X1 U33259 ( .A(n28788), .ZN(p_wishbone_bd_ram_n23542) );
  INV_X1 U33260 ( .A(n61834), .ZN(n28790) );
  INV_X1 U33261 ( .A(n28790), .ZN(p_wishbone_bd_ram_n23541) );
  INV_X1 U33262 ( .A(n61833), .ZN(n28792) );
  INV_X1 U33263 ( .A(n28792), .ZN(p_wishbone_bd_ram_n23540) );
  INV_X1 U33264 ( .A(n61832), .ZN(n28794) );
  INV_X1 U33265 ( .A(n28794), .ZN(p_wishbone_bd_ram_n23539) );
  INV_X1 U33266 ( .A(n61831), .ZN(n28796) );
  INV_X1 U33267 ( .A(n28796), .ZN(p_wishbone_bd_ram_n23538) );
  INV_X1 U33268 ( .A(n61830), .ZN(n28798) );
  INV_X1 U33269 ( .A(n28798), .ZN(p_wishbone_bd_ram_n23537) );
  INV_X1 U33270 ( .A(n61829), .ZN(n28800) );
  INV_X1 U33271 ( .A(n28800), .ZN(p_wishbone_bd_ram_n23536) );
  INV_X1 U33272 ( .A(n61828), .ZN(n28802) );
  INV_X1 U33273 ( .A(n28802), .ZN(p_wishbone_bd_ram_n23535) );
  INV_X1 U33274 ( .A(n61827), .ZN(n28804) );
  INV_X1 U33275 ( .A(n28804), .ZN(p_wishbone_bd_ram_n23534) );
  INV_X1 U33276 ( .A(n61826), .ZN(n28806) );
  INV_X1 U33277 ( .A(n28806), .ZN(p_wishbone_bd_ram_n23533) );
  INV_X1 U33278 ( .A(n61825), .ZN(n28808) );
  INV_X1 U33279 ( .A(n28808), .ZN(p_wishbone_bd_ram_n23532) );
  INV_X1 U33280 ( .A(n61824), .ZN(n28810) );
  INV_X1 U33281 ( .A(n28810), .ZN(p_wishbone_bd_ram_n23531) );
  INV_X1 U33282 ( .A(n61823), .ZN(n28812) );
  INV_X1 U33283 ( .A(n28812), .ZN(p_wishbone_bd_ram_n23530) );
  INV_X1 U33284 ( .A(n61822), .ZN(n28814) );
  INV_X1 U33285 ( .A(n28814), .ZN(p_wishbone_bd_ram_n23529) );
  INV_X1 U33286 ( .A(n61821), .ZN(n28816) );
  INV_X1 U33287 ( .A(n28816), .ZN(p_wishbone_bd_ram_n23528) );
  INV_X1 U33288 ( .A(n61820), .ZN(n28818) );
  INV_X1 U33289 ( .A(n28818), .ZN(p_wishbone_bd_ram_n23527) );
  INV_X1 U33290 ( .A(n61819), .ZN(n28820) );
  INV_X1 U33291 ( .A(n28820), .ZN(p_wishbone_bd_ram_n23526) );
  INV_X1 U33292 ( .A(n61818), .ZN(n28822) );
  INV_X1 U33293 ( .A(n28822), .ZN(p_wishbone_bd_ram_n23525) );
  INV_X1 U33294 ( .A(n61817), .ZN(n28824) );
  INV_X1 U33295 ( .A(n28824), .ZN(p_wishbone_bd_ram_n23524) );
  INV_X1 U33296 ( .A(n61816), .ZN(n28826) );
  INV_X1 U33297 ( .A(n28826), .ZN(p_wishbone_bd_ram_n23523) );
  INV_X1 U33298 ( .A(n61815), .ZN(n28828) );
  INV_X1 U33299 ( .A(n28828), .ZN(p_wishbone_bd_ram_n23522) );
  INV_X1 U33300 ( .A(n61814), .ZN(n28830) );
  INV_X1 U33301 ( .A(n28830), .ZN(p_wishbone_bd_ram_n23521) );
  INV_X1 U33302 ( .A(n61813), .ZN(n28832) );
  INV_X1 U33303 ( .A(n28832), .ZN(p_wishbone_bd_ram_n23520) );
  INV_X1 U33304 ( .A(n61812), .ZN(n28834) );
  INV_X1 U33305 ( .A(n28834), .ZN(p_wishbone_bd_ram_n23519) );
  INV_X1 U33306 ( .A(n61811), .ZN(n28836) );
  INV_X1 U33307 ( .A(n28836), .ZN(p_wishbone_bd_ram_n23518) );
  INV_X1 U33308 ( .A(n61810), .ZN(n28838) );
  INV_X1 U33309 ( .A(n28838), .ZN(p_wishbone_bd_ram_n23517) );
  INV_X1 U33310 ( .A(n61809), .ZN(n28840) );
  INV_X1 U33311 ( .A(n28840), .ZN(p_wishbone_bd_ram_n23516) );
  INV_X1 U33312 ( .A(n61808), .ZN(n28842) );
  INV_X1 U33313 ( .A(n28842), .ZN(p_wishbone_bd_ram_n23515) );
  INV_X1 U33314 ( .A(n61807), .ZN(n28844) );
  INV_X1 U33315 ( .A(n28844), .ZN(p_wishbone_bd_ram_n23514) );
  INV_X1 U33316 ( .A(n61806), .ZN(n28846) );
  INV_X1 U33317 ( .A(n28846), .ZN(p_wishbone_bd_ram_n23513) );
  INV_X1 U33318 ( .A(n61805), .ZN(n28848) );
  INV_X1 U33319 ( .A(n28848), .ZN(p_wishbone_bd_ram_n23512) );
  INV_X1 U33320 ( .A(n61804), .ZN(n28850) );
  INV_X1 U33321 ( .A(n28850), .ZN(p_wishbone_bd_ram_n23511) );
  INV_X1 U33322 ( .A(n61803), .ZN(n28852) );
  INV_X1 U33323 ( .A(n28852), .ZN(p_wishbone_bd_ram_n23510) );
  INV_X1 U33324 ( .A(n61802), .ZN(n28854) );
  INV_X1 U33325 ( .A(n28854), .ZN(p_wishbone_bd_ram_n23509) );
  INV_X1 U33326 ( .A(n61801), .ZN(n28856) );
  INV_X1 U33327 ( .A(n28856), .ZN(p_wishbone_bd_ram_n23508) );
  INV_X1 U33328 ( .A(n61800), .ZN(n28858) );
  INV_X1 U33329 ( .A(n28858), .ZN(p_wishbone_bd_ram_n23507) );
  INV_X1 U33330 ( .A(n61799), .ZN(n28860) );
  INV_X1 U33331 ( .A(n28860), .ZN(p_wishbone_bd_ram_n23506) );
  INV_X1 U33332 ( .A(n61798), .ZN(n28862) );
  INV_X1 U33333 ( .A(n28862), .ZN(p_wishbone_bd_ram_n23505) );
  INV_X1 U33334 ( .A(n61797), .ZN(n28864) );
  INV_X1 U33335 ( .A(n28864), .ZN(p_wishbone_bd_ram_n23504) );
  INV_X1 U33336 ( .A(n61796), .ZN(n28866) );
  INV_X1 U33337 ( .A(n28866), .ZN(p_wishbone_bd_ram_n23503) );
  INV_X1 U33338 ( .A(n61795), .ZN(n28868) );
  INV_X1 U33339 ( .A(n28868), .ZN(p_wishbone_bd_ram_n23502) );
  INV_X1 U33340 ( .A(n61794), .ZN(n28870) );
  INV_X1 U33341 ( .A(n28870), .ZN(p_wishbone_bd_ram_n23501) );
  INV_X1 U33342 ( .A(n61793), .ZN(n28872) );
  INV_X1 U33343 ( .A(n28872), .ZN(p_wishbone_bd_ram_n23500) );
  INV_X1 U33344 ( .A(n61792), .ZN(n28874) );
  INV_X1 U33345 ( .A(n28874), .ZN(p_wishbone_bd_ram_n23499) );
  INV_X1 U33346 ( .A(n61791), .ZN(n28876) );
  INV_X1 U33347 ( .A(n28876), .ZN(p_wishbone_bd_ram_n23498) );
  INV_X1 U33348 ( .A(n61790), .ZN(n28878) );
  INV_X1 U33349 ( .A(n28878), .ZN(p_wishbone_bd_ram_n23497) );
  INV_X1 U33350 ( .A(n61789), .ZN(n28880) );
  INV_X1 U33351 ( .A(n28880), .ZN(p_wishbone_bd_ram_n23496) );
  INV_X1 U33352 ( .A(n61788), .ZN(n28882) );
  INV_X1 U33353 ( .A(n28882), .ZN(p_wishbone_bd_ram_n23495) );
  INV_X1 U33354 ( .A(n61787), .ZN(n28884) );
  INV_X1 U33355 ( .A(n28884), .ZN(p_wishbone_bd_ram_n23494) );
  INV_X1 U33356 ( .A(n61786), .ZN(n28886) );
  INV_X1 U33357 ( .A(n28886), .ZN(p_wishbone_bd_ram_n23493) );
  INV_X1 U33358 ( .A(n61785), .ZN(n28888) );
  INV_X1 U33359 ( .A(n28888), .ZN(p_wishbone_bd_ram_n23492) );
  INV_X1 U33360 ( .A(n61784), .ZN(n28890) );
  INV_X1 U33361 ( .A(n28890), .ZN(p_wishbone_bd_ram_n23491) );
  INV_X1 U33362 ( .A(n61783), .ZN(n28892) );
  INV_X1 U33363 ( .A(n28892), .ZN(p_wishbone_bd_ram_n23490) );
  INV_X1 U33364 ( .A(n61782), .ZN(n28894) );
  INV_X1 U33365 ( .A(n28894), .ZN(p_wishbone_bd_ram_n23489) );
  INV_X1 U33366 ( .A(n61781), .ZN(n28896) );
  INV_X1 U33367 ( .A(n28896), .ZN(p_wishbone_bd_ram_n23488) );
  INV_X1 U33368 ( .A(n61780), .ZN(n28898) );
  INV_X1 U33369 ( .A(n28898), .ZN(p_wishbone_bd_ram_n23487) );
  INV_X1 U33370 ( .A(n61779), .ZN(n28900) );
  INV_X1 U33371 ( .A(n28900), .ZN(p_wishbone_bd_ram_n23486) );
  INV_X1 U33372 ( .A(n61778), .ZN(n28902) );
  INV_X1 U33373 ( .A(n28902), .ZN(p_wishbone_bd_ram_n23485) );
  INV_X1 U33374 ( .A(n61777), .ZN(n28904) );
  INV_X1 U33375 ( .A(n28904), .ZN(p_wishbone_bd_ram_n23484) );
  INV_X1 U33376 ( .A(n61776), .ZN(n28906) );
  INV_X1 U33377 ( .A(n28906), .ZN(p_wishbone_bd_ram_n23483) );
  INV_X1 U33378 ( .A(n61775), .ZN(n28908) );
  INV_X1 U33379 ( .A(n28908), .ZN(p_wishbone_bd_ram_n23482) );
  INV_X1 U33380 ( .A(n61774), .ZN(n28910) );
  INV_X1 U33381 ( .A(n28910), .ZN(p_wishbone_bd_ram_n23481) );
  INV_X1 U33382 ( .A(n61773), .ZN(n28912) );
  INV_X1 U33383 ( .A(n28912), .ZN(p_wishbone_bd_ram_n23480) );
  INV_X1 U33384 ( .A(n61772), .ZN(n28914) );
  INV_X1 U33385 ( .A(n28914), .ZN(p_wishbone_bd_ram_n23479) );
  INV_X1 U33386 ( .A(n61771), .ZN(n28916) );
  INV_X1 U33387 ( .A(n28916), .ZN(p_wishbone_bd_ram_n23478) );
  INV_X1 U33388 ( .A(n61770), .ZN(n28918) );
  INV_X1 U33389 ( .A(n28918), .ZN(p_wishbone_bd_ram_n23477) );
  INV_X1 U33390 ( .A(n61769), .ZN(n28920) );
  INV_X1 U33391 ( .A(n28920), .ZN(p_wishbone_bd_ram_n23476) );
  INV_X1 U33392 ( .A(n61768), .ZN(n28922) );
  INV_X1 U33393 ( .A(n28922), .ZN(p_wishbone_bd_ram_n23475) );
  INV_X1 U33394 ( .A(n61767), .ZN(n28924) );
  INV_X1 U33395 ( .A(n28924), .ZN(p_wishbone_bd_ram_n23474) );
  INV_X1 U33396 ( .A(n61766), .ZN(n28926) );
  INV_X1 U33397 ( .A(n28926), .ZN(p_wishbone_bd_ram_n23473) );
  INV_X1 U33398 ( .A(n61765), .ZN(n28928) );
  INV_X1 U33399 ( .A(n28928), .ZN(p_wishbone_bd_ram_n23472) );
  INV_X1 U33400 ( .A(n61764), .ZN(n28930) );
  INV_X1 U33401 ( .A(n28930), .ZN(p_wishbone_bd_ram_n23471) );
  INV_X1 U33402 ( .A(n61763), .ZN(n28932) );
  INV_X1 U33403 ( .A(n28932), .ZN(p_wishbone_bd_ram_n23470) );
  INV_X1 U33404 ( .A(n61762), .ZN(n28934) );
  INV_X1 U33405 ( .A(n28934), .ZN(p_wishbone_bd_ram_n23469) );
  INV_X1 U33406 ( .A(n61761), .ZN(n28936) );
  INV_X1 U33407 ( .A(n28936), .ZN(p_wishbone_bd_ram_n23468) );
  INV_X1 U33408 ( .A(n61760), .ZN(n28938) );
  INV_X1 U33409 ( .A(n28938), .ZN(p_wishbone_bd_ram_n23467) );
  INV_X1 U33410 ( .A(n61759), .ZN(n28940) );
  INV_X1 U33411 ( .A(n28940), .ZN(p_wishbone_bd_ram_n23466) );
  INV_X1 U33412 ( .A(n61758), .ZN(n28942) );
  INV_X1 U33413 ( .A(n28942), .ZN(p_wishbone_bd_ram_n23465) );
  INV_X1 U33414 ( .A(n61757), .ZN(n28944) );
  INV_X1 U33415 ( .A(n28944), .ZN(p_wishbone_bd_ram_n23464) );
  INV_X1 U33416 ( .A(n61756), .ZN(n28946) );
  INV_X1 U33417 ( .A(n28946), .ZN(p_wishbone_bd_ram_n23463) );
  INV_X1 U33418 ( .A(n61755), .ZN(n28948) );
  INV_X1 U33419 ( .A(n28948), .ZN(p_wishbone_bd_ram_n23462) );
  INV_X1 U33420 ( .A(n61754), .ZN(n28950) );
  INV_X1 U33421 ( .A(n28950), .ZN(p_wishbone_bd_ram_n23461) );
  INV_X1 U33422 ( .A(n61753), .ZN(n28952) );
  INV_X1 U33423 ( .A(n28952), .ZN(p_wishbone_bd_ram_n23460) );
  INV_X1 U33424 ( .A(n61752), .ZN(n28954) );
  INV_X1 U33425 ( .A(n28954), .ZN(p_wishbone_bd_ram_n23459) );
  INV_X1 U33426 ( .A(n61751), .ZN(n28956) );
  INV_X1 U33427 ( .A(n28956), .ZN(p_wishbone_bd_ram_n23458) );
  INV_X1 U33428 ( .A(n61750), .ZN(n28958) );
  INV_X1 U33429 ( .A(n28958), .ZN(p_wishbone_bd_ram_n23457) );
  INV_X1 U33430 ( .A(n61749), .ZN(n28960) );
  INV_X1 U33431 ( .A(n28960), .ZN(p_wishbone_bd_ram_n23456) );
  INV_X1 U33432 ( .A(n61748), .ZN(n28962) );
  INV_X1 U33433 ( .A(n28962), .ZN(p_wishbone_bd_ram_n23455) );
  INV_X1 U33434 ( .A(n61747), .ZN(n28964) );
  INV_X1 U33435 ( .A(n28964), .ZN(p_wishbone_bd_ram_n23454) );
  INV_X1 U33436 ( .A(n61746), .ZN(n28966) );
  INV_X1 U33437 ( .A(n28966), .ZN(p_wishbone_bd_ram_n23453) );
  INV_X1 U33438 ( .A(n61745), .ZN(n28968) );
  INV_X1 U33439 ( .A(n28968), .ZN(p_wishbone_bd_ram_n23452) );
  INV_X1 U33440 ( .A(n61744), .ZN(n28970) );
  INV_X1 U33441 ( .A(n28970), .ZN(p_wishbone_bd_ram_n23451) );
  INV_X1 U33442 ( .A(n61743), .ZN(n28972) );
  INV_X1 U33443 ( .A(n28972), .ZN(p_wishbone_bd_ram_n23450) );
  INV_X1 U33444 ( .A(n61742), .ZN(n28974) );
  INV_X1 U33445 ( .A(n28974), .ZN(p_wishbone_bd_ram_n23449) );
  INV_X1 U33446 ( .A(n61741), .ZN(n28976) );
  INV_X1 U33447 ( .A(n28976), .ZN(p_wishbone_bd_ram_n23448) );
  INV_X1 U33448 ( .A(n61740), .ZN(n28978) );
  INV_X1 U33449 ( .A(n28978), .ZN(p_wishbone_bd_ram_n23447) );
  INV_X1 U33450 ( .A(n61739), .ZN(n28980) );
  INV_X1 U33451 ( .A(n28980), .ZN(p_wishbone_bd_ram_n23446) );
  INV_X1 U33452 ( .A(n61738), .ZN(n28982) );
  INV_X1 U33453 ( .A(n28982), .ZN(p_wishbone_bd_ram_n23445) );
  INV_X1 U33454 ( .A(n61737), .ZN(n28984) );
  INV_X1 U33455 ( .A(n28984), .ZN(p_wishbone_bd_ram_n23444) );
  INV_X1 U33456 ( .A(n61736), .ZN(n28986) );
  INV_X1 U33457 ( .A(n28986), .ZN(p_wishbone_bd_ram_n23443) );
  INV_X1 U33458 ( .A(n61735), .ZN(n28988) );
  INV_X1 U33459 ( .A(n28988), .ZN(p_wishbone_bd_ram_n23442) );
  INV_X1 U33460 ( .A(n61734), .ZN(n28990) );
  INV_X1 U33461 ( .A(n28990), .ZN(p_wishbone_bd_ram_n23441) );
  INV_X1 U33462 ( .A(n61733), .ZN(n28992) );
  INV_X1 U33463 ( .A(n28992), .ZN(p_wishbone_bd_ram_n23440) );
  INV_X1 U33464 ( .A(n61732), .ZN(n28994) );
  INV_X1 U33465 ( .A(n28994), .ZN(p_wishbone_bd_ram_n23439) );
  INV_X1 U33466 ( .A(n61731), .ZN(n28996) );
  INV_X1 U33467 ( .A(n28996), .ZN(p_wishbone_bd_ram_n23438) );
  INV_X1 U33468 ( .A(n61730), .ZN(n28998) );
  INV_X1 U33469 ( .A(n28998), .ZN(p_wishbone_bd_ram_n23437) );
  INV_X1 U33470 ( .A(n61729), .ZN(n29000) );
  INV_X1 U33471 ( .A(n29000), .ZN(p_wishbone_bd_ram_n23436) );
  INV_X1 U33472 ( .A(n61728), .ZN(n29002) );
  INV_X1 U33473 ( .A(n29002), .ZN(p_wishbone_bd_ram_n23435) );
  INV_X1 U33474 ( .A(n61727), .ZN(n29004) );
  INV_X1 U33475 ( .A(n29004), .ZN(p_wishbone_bd_ram_n23434) );
  INV_X1 U33476 ( .A(n61726), .ZN(n29006) );
  INV_X1 U33477 ( .A(n29006), .ZN(p_wishbone_bd_ram_n23433) );
  INV_X1 U33478 ( .A(n61725), .ZN(n29008) );
  INV_X1 U33479 ( .A(n29008), .ZN(p_wishbone_bd_ram_n23432) );
  INV_X1 U33480 ( .A(n61724), .ZN(n29010) );
  INV_X1 U33481 ( .A(n29010), .ZN(p_wishbone_bd_ram_n23431) );
  INV_X1 U33482 ( .A(n61723), .ZN(n29012) );
  INV_X1 U33483 ( .A(n29012), .ZN(p_wishbone_bd_ram_n23430) );
  INV_X1 U33484 ( .A(n61722), .ZN(n29014) );
  INV_X1 U33485 ( .A(n29014), .ZN(p_wishbone_bd_ram_n23429) );
  INV_X1 U33486 ( .A(n61721), .ZN(n29016) );
  INV_X1 U33487 ( .A(n29016), .ZN(p_wishbone_bd_ram_n23428) );
  INV_X1 U33488 ( .A(n61720), .ZN(n29018) );
  INV_X1 U33489 ( .A(n29018), .ZN(p_wishbone_bd_ram_n23427) );
  INV_X1 U33490 ( .A(n61719), .ZN(n29020) );
  INV_X1 U33491 ( .A(n29020), .ZN(p_wishbone_bd_ram_n23426) );
  INV_X1 U33492 ( .A(n61718), .ZN(n29022) );
  INV_X1 U33493 ( .A(n29022), .ZN(p_wishbone_bd_ram_n23425) );
  INV_X1 U33494 ( .A(n61717), .ZN(n29024) );
  INV_X1 U33495 ( .A(n29024), .ZN(p_wishbone_bd_ram_n23424) );
  INV_X1 U33496 ( .A(n61716), .ZN(n29026) );
  INV_X1 U33497 ( .A(n29026), .ZN(p_wishbone_bd_ram_n23423) );
  INV_X1 U33498 ( .A(n61715), .ZN(n29028) );
  INV_X1 U33499 ( .A(n29028), .ZN(p_wishbone_bd_ram_n23422) );
  INV_X1 U33500 ( .A(n61714), .ZN(n29030) );
  INV_X1 U33501 ( .A(n29030), .ZN(p_wishbone_bd_ram_n23421) );
  INV_X1 U33502 ( .A(n61713), .ZN(n29032) );
  INV_X1 U33503 ( .A(n29032), .ZN(p_wishbone_bd_ram_n23420) );
  INV_X1 U33504 ( .A(n61712), .ZN(n29034) );
  INV_X1 U33505 ( .A(n29034), .ZN(p_wishbone_bd_ram_n23419) );
  INV_X1 U33506 ( .A(n61711), .ZN(n29036) );
  INV_X1 U33507 ( .A(n29036), .ZN(p_wishbone_bd_ram_n23418) );
  INV_X1 U33508 ( .A(n61710), .ZN(n29038) );
  INV_X1 U33509 ( .A(n29038), .ZN(p_wishbone_bd_ram_n23417) );
  INV_X1 U33510 ( .A(n61709), .ZN(n29040) );
  INV_X1 U33511 ( .A(n29040), .ZN(p_wishbone_bd_ram_n23416) );
  INV_X1 U33512 ( .A(n61708), .ZN(n29042) );
  INV_X1 U33513 ( .A(n29042), .ZN(p_wishbone_bd_ram_n23415) );
  INV_X1 U33514 ( .A(n61707), .ZN(n29044) );
  INV_X1 U33515 ( .A(n29044), .ZN(p_wishbone_bd_ram_n23414) );
  INV_X1 U33516 ( .A(n61706), .ZN(n29046) );
  INV_X1 U33517 ( .A(n29046), .ZN(p_wishbone_bd_ram_n23413) );
  INV_X1 U33518 ( .A(n61705), .ZN(n29048) );
  INV_X1 U33519 ( .A(n29048), .ZN(p_wishbone_bd_ram_n23412) );
  INV_X1 U33520 ( .A(n61704), .ZN(n29050) );
  INV_X1 U33521 ( .A(n29050), .ZN(p_wishbone_bd_ram_n23411) );
  INV_X1 U33522 ( .A(n61703), .ZN(n29052) );
  INV_X1 U33523 ( .A(n29052), .ZN(p_wishbone_bd_ram_n23410) );
  INV_X1 U33524 ( .A(n61702), .ZN(n29054) );
  INV_X1 U33525 ( .A(n29054), .ZN(p_wishbone_bd_ram_n23409) );
  INV_X1 U33526 ( .A(n61701), .ZN(n29056) );
  INV_X1 U33527 ( .A(n29056), .ZN(p_wishbone_bd_ram_n23408) );
  INV_X1 U33528 ( .A(n61700), .ZN(n29058) );
  INV_X1 U33529 ( .A(n29058), .ZN(p_wishbone_bd_ram_n23407) );
  INV_X1 U33530 ( .A(n61699), .ZN(n29060) );
  INV_X1 U33531 ( .A(n29060), .ZN(p_wishbone_bd_ram_n23406) );
  INV_X1 U33532 ( .A(n61698), .ZN(n29062) );
  INV_X1 U33533 ( .A(n29062), .ZN(p_wishbone_bd_ram_n23405) );
  INV_X1 U33534 ( .A(n61697), .ZN(n29064) );
  INV_X1 U33535 ( .A(n29064), .ZN(p_wishbone_bd_ram_n23404) );
  INV_X1 U33536 ( .A(n61696), .ZN(n29066) );
  INV_X1 U33537 ( .A(n29066), .ZN(p_wishbone_bd_ram_n23403) );
  INV_X1 U33538 ( .A(n61695), .ZN(n29068) );
  INV_X1 U33539 ( .A(n29068), .ZN(p_wishbone_bd_ram_n23402) );
  INV_X1 U33540 ( .A(n61694), .ZN(n29070) );
  INV_X1 U33541 ( .A(n29070), .ZN(p_wishbone_bd_ram_n23401) );
  INV_X1 U33542 ( .A(n61693), .ZN(n29072) );
  INV_X1 U33543 ( .A(n29072), .ZN(p_wishbone_bd_ram_n23400) );
  INV_X1 U33544 ( .A(n61692), .ZN(n29074) );
  INV_X1 U33545 ( .A(n29074), .ZN(p_wishbone_bd_ram_n23399) );
  INV_X1 U33546 ( .A(n61691), .ZN(n29076) );
  INV_X1 U33547 ( .A(n29076), .ZN(p_wishbone_bd_ram_n23398) );
  INV_X1 U33548 ( .A(n61690), .ZN(n29078) );
  INV_X1 U33549 ( .A(n29078), .ZN(p_wishbone_bd_ram_n23397) );
  INV_X1 U33550 ( .A(n61689), .ZN(n29080) );
  INV_X1 U33551 ( .A(n29080), .ZN(p_wishbone_bd_ram_n23396) );
  INV_X1 U33552 ( .A(n61688), .ZN(n29082) );
  INV_X1 U33553 ( .A(n29082), .ZN(p_wishbone_bd_ram_n23395) );
  INV_X1 U33554 ( .A(n61687), .ZN(n29084) );
  INV_X1 U33555 ( .A(n29084), .ZN(p_wishbone_bd_ram_n23394) );
  INV_X1 U33556 ( .A(n61686), .ZN(n29086) );
  INV_X1 U33557 ( .A(n29086), .ZN(p_wishbone_bd_ram_n23393) );
  INV_X1 U33558 ( .A(n61685), .ZN(n29088) );
  INV_X1 U33559 ( .A(n29088), .ZN(p_wishbone_bd_ram_n23392) );
  INV_X1 U33560 ( .A(n61684), .ZN(n29090) );
  INV_X1 U33561 ( .A(n29090), .ZN(p_wishbone_bd_ram_n23391) );
  INV_X1 U33562 ( .A(n61683), .ZN(n29092) );
  INV_X1 U33563 ( .A(n29092), .ZN(p_wishbone_bd_ram_n23390) );
  INV_X1 U33564 ( .A(n61682), .ZN(n29094) );
  INV_X1 U33565 ( .A(n29094), .ZN(p_wishbone_bd_ram_n23389) );
  INV_X1 U33566 ( .A(n61681), .ZN(n29096) );
  INV_X1 U33567 ( .A(n29096), .ZN(p_wishbone_bd_ram_n23388) );
  INV_X1 U33568 ( .A(n61680), .ZN(n29098) );
  INV_X1 U33569 ( .A(n29098), .ZN(p_wishbone_bd_ram_n23387) );
  INV_X1 U33570 ( .A(n61679), .ZN(n29100) );
  INV_X1 U33571 ( .A(n29100), .ZN(p_wishbone_bd_ram_n23386) );
  INV_X1 U33572 ( .A(n61678), .ZN(n29102) );
  INV_X1 U33573 ( .A(n29102), .ZN(p_wishbone_bd_ram_n23385) );
  INV_X1 U33574 ( .A(n61677), .ZN(n29104) );
  INV_X1 U33575 ( .A(n29104), .ZN(p_wishbone_bd_ram_n23384) );
  INV_X1 U33576 ( .A(n61676), .ZN(n29106) );
  INV_X1 U33577 ( .A(n29106), .ZN(p_wishbone_bd_ram_n23383) );
  INV_X1 U33578 ( .A(n61675), .ZN(n29108) );
  INV_X1 U33579 ( .A(n29108), .ZN(p_wishbone_bd_ram_n23382) );
  INV_X1 U33580 ( .A(n61674), .ZN(n29110) );
  INV_X1 U33581 ( .A(n29110), .ZN(p_wishbone_bd_ram_n23381) );
  INV_X1 U33582 ( .A(n61673), .ZN(n29112) );
  INV_X1 U33583 ( .A(n29112), .ZN(p_wishbone_bd_ram_n23380) );
  INV_X1 U33584 ( .A(n61672), .ZN(n29114) );
  INV_X1 U33585 ( .A(n29114), .ZN(p_wishbone_bd_ram_n23379) );
  INV_X1 U33586 ( .A(n61671), .ZN(n29116) );
  INV_X1 U33587 ( .A(n29116), .ZN(p_wishbone_bd_ram_n23378) );
  INV_X1 U33588 ( .A(n61670), .ZN(n29118) );
  INV_X1 U33589 ( .A(n29118), .ZN(p_wishbone_bd_ram_n23377) );
  INV_X1 U33590 ( .A(n61669), .ZN(n29120) );
  INV_X1 U33591 ( .A(n29120), .ZN(p_wishbone_bd_ram_n23376) );
  INV_X1 U33592 ( .A(n61668), .ZN(n29122) );
  INV_X1 U33593 ( .A(n29122), .ZN(p_wishbone_bd_ram_n23375) );
  INV_X1 U33594 ( .A(n61667), .ZN(n29124) );
  INV_X1 U33595 ( .A(n29124), .ZN(p_wishbone_bd_ram_n23374) );
  INV_X1 U33596 ( .A(n61666), .ZN(n29126) );
  INV_X1 U33597 ( .A(n29126), .ZN(p_wishbone_bd_ram_n23373) );
  INV_X1 U33598 ( .A(n61665), .ZN(n29128) );
  INV_X1 U33599 ( .A(n29128), .ZN(p_wishbone_bd_ram_n23372) );
  INV_X1 U33600 ( .A(n61664), .ZN(n29130) );
  INV_X1 U33601 ( .A(n29130), .ZN(p_wishbone_bd_ram_n23371) );
  INV_X1 U33602 ( .A(n61663), .ZN(n29132) );
  INV_X1 U33603 ( .A(n29132), .ZN(p_wishbone_bd_ram_n23370) );
  INV_X1 U33604 ( .A(n61662), .ZN(n29134) );
  INV_X1 U33605 ( .A(n29134), .ZN(p_wishbone_bd_ram_n23369) );
  INV_X1 U33606 ( .A(n61661), .ZN(n29136) );
  INV_X1 U33607 ( .A(n29136), .ZN(p_wishbone_bd_ram_n23368) );
  INV_X1 U33608 ( .A(n61660), .ZN(n29138) );
  INV_X1 U33609 ( .A(n29138), .ZN(p_wishbone_bd_ram_n23367) );
  INV_X1 U33610 ( .A(n61659), .ZN(n29140) );
  INV_X1 U33611 ( .A(n29140), .ZN(p_wishbone_bd_ram_n23366) );
  INV_X1 U33612 ( .A(n61658), .ZN(n29142) );
  INV_X1 U33613 ( .A(n29142), .ZN(p_wishbone_bd_ram_n23365) );
  INV_X1 U33614 ( .A(n61657), .ZN(n29144) );
  INV_X1 U33615 ( .A(n29144), .ZN(p_wishbone_bd_ram_n23364) );
  INV_X1 U33616 ( .A(n61656), .ZN(n29146) );
  INV_X1 U33617 ( .A(n29146), .ZN(p_wishbone_bd_ram_n23363) );
  INV_X1 U33618 ( .A(n61655), .ZN(n29148) );
  INV_X1 U33619 ( .A(n29148), .ZN(p_wishbone_bd_ram_n23362) );
  INV_X1 U33620 ( .A(n61654), .ZN(n29150) );
  INV_X1 U33621 ( .A(n29150), .ZN(p_wishbone_bd_ram_n23361) );
  INV_X1 U33622 ( .A(n61653), .ZN(n29152) );
  INV_X1 U33623 ( .A(n29152), .ZN(p_wishbone_bd_ram_n23360) );
  INV_X1 U33624 ( .A(n61652), .ZN(n29154) );
  INV_X1 U33625 ( .A(n29154), .ZN(p_wishbone_bd_ram_n23359) );
  INV_X1 U33626 ( .A(n61651), .ZN(n29156) );
  INV_X1 U33627 ( .A(n29156), .ZN(p_wishbone_bd_ram_n23358) );
  INV_X1 U33628 ( .A(n61650), .ZN(n29158) );
  INV_X1 U33629 ( .A(n29158), .ZN(p_wishbone_bd_ram_n23357) );
  INV_X1 U33630 ( .A(n61649), .ZN(n29160) );
  INV_X1 U33631 ( .A(n29160), .ZN(p_wishbone_bd_ram_n23356) );
  INV_X1 U33632 ( .A(n61648), .ZN(n29162) );
  INV_X1 U33633 ( .A(n29162), .ZN(p_wishbone_bd_ram_n23355) );
  INV_X1 U33634 ( .A(n61647), .ZN(n29164) );
  INV_X1 U33635 ( .A(n29164), .ZN(p_wishbone_bd_ram_n23354) );
  INV_X1 U33636 ( .A(n61646), .ZN(n29166) );
  INV_X1 U33637 ( .A(n29166), .ZN(p_wishbone_bd_ram_n23353) );
  INV_X1 U33638 ( .A(n61645), .ZN(n29168) );
  INV_X1 U33639 ( .A(n29168), .ZN(p_wishbone_bd_ram_n23352) );
  INV_X1 U33640 ( .A(n61644), .ZN(n29170) );
  INV_X1 U33641 ( .A(n29170), .ZN(p_wishbone_bd_ram_n23351) );
  INV_X1 U33642 ( .A(n61643), .ZN(n29172) );
  INV_X1 U33643 ( .A(n29172), .ZN(p_wishbone_bd_ram_n23350) );
  INV_X1 U33644 ( .A(n61642), .ZN(n29174) );
  INV_X1 U33645 ( .A(n29174), .ZN(p_wishbone_bd_ram_n23349) );
  INV_X1 U33646 ( .A(n61641), .ZN(n29176) );
  INV_X1 U33647 ( .A(n29176), .ZN(p_wishbone_bd_ram_n23348) );
  INV_X1 U33648 ( .A(n61640), .ZN(n29178) );
  INV_X1 U33649 ( .A(n29178), .ZN(p_wishbone_bd_ram_n23347) );
  INV_X1 U33650 ( .A(n61639), .ZN(n29180) );
  INV_X1 U33651 ( .A(n29180), .ZN(p_wishbone_bd_ram_n23346) );
  INV_X1 U33652 ( .A(n61638), .ZN(n29182) );
  INV_X1 U33653 ( .A(n29182), .ZN(p_wishbone_bd_ram_n23345) );
  INV_X1 U33654 ( .A(n61637), .ZN(n29184) );
  INV_X1 U33655 ( .A(n29184), .ZN(p_wishbone_bd_ram_n23344) );
  INV_X1 U33656 ( .A(n61636), .ZN(n29186) );
  INV_X1 U33657 ( .A(n29186), .ZN(p_wishbone_bd_ram_n23343) );
  INV_X1 U33658 ( .A(n61635), .ZN(n29188) );
  INV_X1 U33659 ( .A(n29188), .ZN(p_wishbone_bd_ram_n23342) );
  INV_X1 U33660 ( .A(n61634), .ZN(n29190) );
  INV_X1 U33661 ( .A(n29190), .ZN(p_wishbone_bd_ram_n23341) );
  INV_X1 U33662 ( .A(n61633), .ZN(n29192) );
  INV_X1 U33663 ( .A(n29192), .ZN(p_wishbone_bd_ram_n23340) );
  INV_X1 U33664 ( .A(n61632), .ZN(n29194) );
  INV_X1 U33665 ( .A(n29194), .ZN(p_wishbone_bd_ram_n23339) );
  INV_X1 U33666 ( .A(n61631), .ZN(n29196) );
  INV_X1 U33667 ( .A(n29196), .ZN(p_wishbone_bd_ram_n23338) );
  INV_X1 U33668 ( .A(n61630), .ZN(n29198) );
  INV_X1 U33669 ( .A(n29198), .ZN(p_wishbone_bd_ram_n23337) );
  INV_X1 U33670 ( .A(n61629), .ZN(n29200) );
  INV_X1 U33671 ( .A(n29200), .ZN(p_wishbone_bd_ram_n23336) );
  INV_X1 U33672 ( .A(n61628), .ZN(n29202) );
  INV_X1 U33673 ( .A(n29202), .ZN(p_wishbone_bd_ram_n23335) );
  INV_X1 U33674 ( .A(n61627), .ZN(n29204) );
  INV_X1 U33675 ( .A(n29204), .ZN(p_wishbone_bd_ram_n23334) );
  INV_X1 U33676 ( .A(n61626), .ZN(n29206) );
  INV_X1 U33677 ( .A(n29206), .ZN(p_wishbone_bd_ram_n23333) );
  INV_X1 U33678 ( .A(n61625), .ZN(n29208) );
  INV_X1 U33679 ( .A(n29208), .ZN(p_wishbone_bd_ram_n23332) );
  INV_X1 U33680 ( .A(n61624), .ZN(n29210) );
  INV_X1 U33681 ( .A(n29210), .ZN(p_wishbone_bd_ram_n23331) );
  INV_X1 U33682 ( .A(n61623), .ZN(n29212) );
  INV_X1 U33683 ( .A(n29212), .ZN(p_wishbone_bd_ram_n23330) );
  INV_X1 U33684 ( .A(n61622), .ZN(n29214) );
  INV_X1 U33685 ( .A(n29214), .ZN(p_wishbone_bd_ram_n23329) );
  INV_X1 U33686 ( .A(n61621), .ZN(n29216) );
  INV_X1 U33687 ( .A(n29216), .ZN(p_wishbone_bd_ram_n23328) );
  INV_X1 U33688 ( .A(n61620), .ZN(n29218) );
  INV_X1 U33689 ( .A(n29218), .ZN(p_wishbone_bd_ram_n23327) );
  INV_X1 U33690 ( .A(n61619), .ZN(n29220) );
  INV_X1 U33691 ( .A(n29220), .ZN(p_wishbone_bd_ram_n23326) );
  INV_X1 U33692 ( .A(n61618), .ZN(n29222) );
  INV_X1 U33693 ( .A(n29222), .ZN(p_wishbone_bd_ram_n23325) );
  INV_X1 U33694 ( .A(n61617), .ZN(n29224) );
  INV_X1 U33695 ( .A(n29224), .ZN(p_wishbone_bd_ram_n23324) );
  INV_X1 U33696 ( .A(n61616), .ZN(n29226) );
  INV_X1 U33697 ( .A(n29226), .ZN(p_wishbone_bd_ram_n23323) );
  INV_X1 U33698 ( .A(n61615), .ZN(n29228) );
  INV_X1 U33699 ( .A(n29228), .ZN(p_wishbone_bd_ram_n23322) );
  INV_X1 U33700 ( .A(n61614), .ZN(n29230) );
  INV_X1 U33701 ( .A(n29230), .ZN(p_wishbone_bd_ram_n23321) );
  INV_X1 U33702 ( .A(n61613), .ZN(n29232) );
  INV_X1 U33703 ( .A(n29232), .ZN(p_wishbone_bd_ram_n23320) );
  INV_X1 U33704 ( .A(n61612), .ZN(n29234) );
  INV_X1 U33705 ( .A(n29234), .ZN(p_wishbone_bd_ram_n23319) );
  INV_X1 U33706 ( .A(n61611), .ZN(n29236) );
  INV_X1 U33707 ( .A(n29236), .ZN(p_wishbone_bd_ram_n23318) );
  INV_X1 U33708 ( .A(n61610), .ZN(n29238) );
  INV_X1 U33709 ( .A(n29238), .ZN(p_wishbone_bd_ram_n23317) );
  INV_X1 U33710 ( .A(n61609), .ZN(n29240) );
  INV_X1 U33711 ( .A(n29240), .ZN(p_wishbone_bd_ram_n23316) );
  INV_X1 U33712 ( .A(n61608), .ZN(n29242) );
  INV_X1 U33713 ( .A(n29242), .ZN(p_wishbone_bd_ram_n23315) );
  INV_X1 U33714 ( .A(n61607), .ZN(n29244) );
  INV_X1 U33715 ( .A(n29244), .ZN(p_wishbone_bd_ram_n23314) );
  INV_X1 U33716 ( .A(n61606), .ZN(n29246) );
  INV_X1 U33717 ( .A(n29246), .ZN(p_wishbone_bd_ram_n23313) );
  INV_X1 U33718 ( .A(n61605), .ZN(n29248) );
  INV_X1 U33719 ( .A(n29248), .ZN(p_wishbone_bd_ram_n23311) );
  INV_X1 U33720 ( .A(n61604), .ZN(n29250) );
  INV_X1 U33721 ( .A(n29250), .ZN(p_wishbone_bd_ram_n23309) );
  INV_X1 U33722 ( .A(n61603), .ZN(n29252) );
  INV_X1 U33723 ( .A(n29252), .ZN(p_wishbone_bd_ram_n23308) );
  INV_X1 U33724 ( .A(n61602), .ZN(n29254) );
  INV_X1 U33725 ( .A(n29254), .ZN(p_wishbone_bd_ram_n23306) );
  INV_X1 U33726 ( .A(n61601), .ZN(n29256) );
  INV_X1 U33727 ( .A(n29256), .ZN(p_wishbone_bd_ram_n23304) );
  INV_X1 U33728 ( .A(n61600), .ZN(n29258) );
  INV_X1 U33729 ( .A(n29258), .ZN(p_wishbone_bd_ram_n23303) );
  INV_X1 U33730 ( .A(n61599), .ZN(n29260) );
  INV_X1 U33731 ( .A(n29260), .ZN(p_wishbone_bd_ram_n23302) );
  INV_X1 U33732 ( .A(n61598), .ZN(n29262) );
  INV_X1 U33733 ( .A(n29262), .ZN(p_wishbone_bd_ram_n23301) );
  INV_X1 U33734 ( .A(n61597), .ZN(n29264) );
  INV_X1 U33735 ( .A(n29264), .ZN(p_wishbone_bd_ram_n23300) );
  INV_X1 U33736 ( .A(n61596), .ZN(n29266) );
  INV_X1 U33737 ( .A(n29266), .ZN(p_wishbone_bd_ram_n23299) );
  INV_X1 U33738 ( .A(n61595), .ZN(n29268) );
  INV_X1 U33739 ( .A(n29268), .ZN(p_wishbone_bd_ram_n23298) );
  INV_X1 U33740 ( .A(n61594), .ZN(n29270) );
  INV_X1 U33741 ( .A(n29270), .ZN(p_wishbone_bd_ram_n23297) );
  INV_X1 U33742 ( .A(n61593), .ZN(n29272) );
  INV_X1 U33743 ( .A(n29272), .ZN(p_wishbone_bd_ram_n23296) );
  INV_X1 U33744 ( .A(n61592), .ZN(n29274) );
  INV_X1 U33745 ( .A(n29274), .ZN(p_wishbone_bd_ram_n23295) );
  INV_X1 U33746 ( .A(n61591), .ZN(n29276) );
  INV_X1 U33747 ( .A(n29276), .ZN(p_wishbone_bd_ram_n23294) );
  INV_X1 U33748 ( .A(n61590), .ZN(n29278) );
  INV_X1 U33749 ( .A(n29278), .ZN(p_wishbone_bd_ram_n23293) );
  INV_X1 U33750 ( .A(n61589), .ZN(n29280) );
  INV_X1 U33751 ( .A(n29280), .ZN(p_wishbone_bd_ram_n23292) );
  INV_X1 U33752 ( .A(n61588), .ZN(n29282) );
  INV_X1 U33753 ( .A(n29282), .ZN(p_wishbone_bd_ram_n23291) );
  INV_X1 U33754 ( .A(n61587), .ZN(n29284) );
  INV_X1 U33755 ( .A(n29284), .ZN(p_wishbone_bd_ram_n23290) );
  INV_X1 U33756 ( .A(n61586), .ZN(n29286) );
  INV_X1 U33757 ( .A(n29286), .ZN(p_wishbone_bd_ram_n23289) );
  INV_X1 U33758 ( .A(n61585), .ZN(n29288) );
  INV_X1 U33759 ( .A(n29288), .ZN(p_wishbone_bd_ram_n23288) );
  INV_X1 U33760 ( .A(n61584), .ZN(n29290) );
  INV_X1 U33761 ( .A(n29290), .ZN(p_wishbone_bd_ram_n23287) );
  INV_X1 U33762 ( .A(n61583), .ZN(n29292) );
  INV_X1 U33763 ( .A(n29292), .ZN(p_wishbone_bd_ram_n23286) );
  INV_X1 U33764 ( .A(n61582), .ZN(n29294) );
  INV_X1 U33765 ( .A(n29294), .ZN(p_wishbone_bd_ram_n23285) );
  INV_X1 U33766 ( .A(n61581), .ZN(n29296) );
  INV_X1 U33767 ( .A(n29296), .ZN(p_wishbone_bd_ram_n23284) );
  INV_X1 U33768 ( .A(n61580), .ZN(n29298) );
  INV_X1 U33769 ( .A(n29298), .ZN(p_wishbone_bd_ram_n23283) );
  INV_X1 U33770 ( .A(n61579), .ZN(n29300) );
  INV_X1 U33771 ( .A(n29300), .ZN(p_wishbone_bd_ram_n23282) );
  INV_X1 U33772 ( .A(n61578), .ZN(n29302) );
  INV_X1 U33773 ( .A(n29302), .ZN(p_wishbone_bd_ram_n23281) );
  INV_X1 U33774 ( .A(n61577), .ZN(n29304) );
  INV_X1 U33775 ( .A(n29304), .ZN(p_wishbone_bd_ram_n23280) );
  INV_X1 U33776 ( .A(n61576), .ZN(n29306) );
  INV_X1 U33777 ( .A(n29306), .ZN(p_wishbone_bd_ram_n23279) );
  INV_X1 U33778 ( .A(n61575), .ZN(n29308) );
  INV_X1 U33779 ( .A(n29308), .ZN(p_wishbone_bd_ram_n23278) );
  INV_X1 U33780 ( .A(n61574), .ZN(n29310) );
  INV_X1 U33781 ( .A(n29310), .ZN(p_wishbone_bd_ram_n23277) );
  INV_X1 U33782 ( .A(n61573), .ZN(n29312) );
  INV_X1 U33783 ( .A(n29312), .ZN(p_wishbone_bd_ram_n23276) );
  INV_X1 U33784 ( .A(n61572), .ZN(n29314) );
  INV_X1 U33785 ( .A(n29314), .ZN(p_wishbone_bd_ram_n23275) );
  INV_X1 U33786 ( .A(n61571), .ZN(n29316) );
  INV_X1 U33787 ( .A(n29316), .ZN(p_wishbone_bd_ram_n23274) );
  INV_X1 U33788 ( .A(n61570), .ZN(n29318) );
  INV_X1 U33789 ( .A(n29318), .ZN(p_wishbone_bd_ram_n23273) );
  INV_X1 U33790 ( .A(n61569), .ZN(n29320) );
  INV_X1 U33791 ( .A(n29320), .ZN(p_wishbone_bd_ram_n23272) );
  INV_X1 U33792 ( .A(n61568), .ZN(n29322) );
  INV_X1 U33793 ( .A(n29322), .ZN(p_wishbone_bd_ram_n23271) );
  INV_X1 U33794 ( .A(n61567), .ZN(n29324) );
  INV_X1 U33795 ( .A(n29324), .ZN(p_wishbone_bd_ram_n23270) );
  INV_X1 U33796 ( .A(n61566), .ZN(n29326) );
  INV_X1 U33797 ( .A(n29326), .ZN(p_wishbone_bd_ram_n23269) );
  INV_X1 U33798 ( .A(n61565), .ZN(n29328) );
  INV_X1 U33799 ( .A(n29328), .ZN(p_wishbone_bd_ram_n23268) );
  INV_X1 U33800 ( .A(n61564), .ZN(n29330) );
  INV_X1 U33801 ( .A(n29330), .ZN(p_wishbone_bd_ram_n23267) );
  INV_X1 U33802 ( .A(n61563), .ZN(n29332) );
  INV_X1 U33803 ( .A(n29332), .ZN(p_wishbone_bd_ram_n23266) );
  INV_X1 U33804 ( .A(n61562), .ZN(n29334) );
  INV_X1 U33805 ( .A(n29334), .ZN(p_wishbone_bd_ram_n23265) );
  INV_X1 U33806 ( .A(n61561), .ZN(n29336) );
  INV_X1 U33807 ( .A(n29336), .ZN(p_wishbone_bd_ram_n23264) );
  INV_X1 U33808 ( .A(n61560), .ZN(n29338) );
  INV_X1 U33809 ( .A(n29338), .ZN(p_wishbone_bd_ram_n23262) );
  INV_X1 U33810 ( .A(n61559), .ZN(n29340) );
  INV_X1 U33811 ( .A(n29340), .ZN(p_wishbone_bd_ram_n23259) );
  INV_X1 U33812 ( .A(n61558), .ZN(n29342) );
  INV_X1 U33813 ( .A(n29342), .ZN(p_wishbone_bd_ram_n23257) );
  INV_X1 U33814 ( .A(n61557), .ZN(n29344) );
  INV_X1 U33815 ( .A(n29344), .ZN(p_wishbone_bd_ram_n23256) );
  INV_X1 U33816 ( .A(n61556), .ZN(n29346) );
  INV_X1 U33817 ( .A(n29346), .ZN(p_wishbone_bd_ram_n23255) );
  INV_X1 U33818 ( .A(n61555), .ZN(n29348) );
  INV_X1 U33819 ( .A(n29348), .ZN(p_wishbone_bd_ram_n23254) );
  INV_X1 U33820 ( .A(n61554), .ZN(n29350) );
  INV_X1 U33821 ( .A(n29350), .ZN(p_wishbone_bd_ram_n23253) );
  INV_X1 U33822 ( .A(n61553), .ZN(n29352) );
  INV_X1 U33823 ( .A(n29352), .ZN(p_wishbone_bd_ram_n23252) );
  INV_X1 U33824 ( .A(n61552), .ZN(n29354) );
  INV_X1 U33825 ( .A(n29354), .ZN(p_wishbone_bd_ram_n23251) );
  INV_X1 U33826 ( .A(n61551), .ZN(n29356) );
  INV_X1 U33827 ( .A(n29356), .ZN(p_wishbone_bd_ram_n23250) );
  INV_X1 U33828 ( .A(n61550), .ZN(n29358) );
  INV_X1 U33829 ( .A(n29358), .ZN(p_wishbone_bd_ram_n23249) );
  INV_X1 U33830 ( .A(n61549), .ZN(n29360) );
  INV_X1 U33831 ( .A(n29360), .ZN(p_wishbone_bd_ram_n23248) );
  INV_X1 U33832 ( .A(n61548), .ZN(n29362) );
  INV_X1 U33833 ( .A(n29362), .ZN(p_wishbone_bd_ram_n23247) );
  INV_X1 U33834 ( .A(n61547), .ZN(n29364) );
  INV_X1 U33835 ( .A(n29364), .ZN(p_wishbone_bd_ram_n23246) );
  INV_X1 U33836 ( .A(n61546), .ZN(n29366) );
  INV_X1 U33837 ( .A(n29366), .ZN(p_wishbone_bd_ram_n23245) );
  INV_X1 U33838 ( .A(n61545), .ZN(n29368) );
  INV_X1 U33839 ( .A(n29368), .ZN(p_wishbone_bd_ram_n23244) );
  INV_X1 U33840 ( .A(n61544), .ZN(n29370) );
  INV_X1 U33841 ( .A(n29370), .ZN(p_wishbone_bd_ram_n23243) );
  INV_X1 U33842 ( .A(n61543), .ZN(n29372) );
  INV_X1 U33843 ( .A(n29372), .ZN(p_wishbone_bd_ram_n23242) );
  INV_X1 U33844 ( .A(n61542), .ZN(n29374) );
  INV_X1 U33845 ( .A(n29374), .ZN(p_wishbone_bd_ram_n23241) );
  INV_X1 U33846 ( .A(n61541), .ZN(n29376) );
  INV_X1 U33847 ( .A(n29376), .ZN(p_wishbone_bd_ram_n23240) );
  INV_X1 U33848 ( .A(n61540), .ZN(n29378) );
  INV_X1 U33849 ( .A(n29378), .ZN(p_wishbone_bd_ram_n23239) );
  INV_X1 U33850 ( .A(n61539), .ZN(n29380) );
  INV_X1 U33851 ( .A(n29380), .ZN(p_wishbone_bd_ram_n23238) );
  INV_X1 U33852 ( .A(n61538), .ZN(n29382) );
  INV_X1 U33853 ( .A(n29382), .ZN(p_wishbone_bd_ram_n23237) );
  INV_X1 U33854 ( .A(n61537), .ZN(n29384) );
  INV_X1 U33855 ( .A(n29384), .ZN(p_wishbone_bd_ram_n23236) );
  INV_X1 U33856 ( .A(n61536), .ZN(n29386) );
  INV_X1 U33857 ( .A(n29386), .ZN(p_wishbone_bd_ram_n23235) );
  INV_X1 U33858 ( .A(n61535), .ZN(n29388) );
  INV_X1 U33859 ( .A(n29388), .ZN(p_wishbone_bd_ram_n23234) );
  INV_X1 U33860 ( .A(n61534), .ZN(n29390) );
  INV_X1 U33861 ( .A(n29390), .ZN(p_wishbone_bd_ram_n23233) );
  INV_X1 U33862 ( .A(n61533), .ZN(n29392) );
  INV_X1 U33863 ( .A(n29392), .ZN(p_wishbone_bd_ram_n23232) );
  INV_X1 U33864 ( .A(n61532), .ZN(n29394) );
  INV_X1 U33865 ( .A(n29394), .ZN(p_wishbone_bd_ram_n23231) );
  INV_X1 U33866 ( .A(n61531), .ZN(n29396) );
  INV_X1 U33867 ( .A(n29396), .ZN(p_wishbone_bd_ram_n23230) );
  INV_X1 U33868 ( .A(n61530), .ZN(n29398) );
  INV_X1 U33869 ( .A(n29398), .ZN(p_wishbone_bd_ram_n23229) );
  INV_X1 U33870 ( .A(n61529), .ZN(n29400) );
  INV_X1 U33871 ( .A(n29400), .ZN(p_wishbone_bd_ram_n23228) );
  INV_X1 U33872 ( .A(n61528), .ZN(n29402) );
  INV_X1 U33873 ( .A(n29402), .ZN(p_wishbone_bd_ram_n23227) );
  INV_X1 U33874 ( .A(n61527), .ZN(n29404) );
  INV_X1 U33875 ( .A(n29404), .ZN(p_wishbone_bd_ram_n23226) );
  INV_X1 U33876 ( .A(n61526), .ZN(n29406) );
  INV_X1 U33877 ( .A(n29406), .ZN(p_wishbone_bd_ram_n23225) );
  INV_X1 U33878 ( .A(n61525), .ZN(n29408) );
  INV_X1 U33879 ( .A(n29408), .ZN(p_wishbone_bd_ram_n23224) );
  INV_X1 U33880 ( .A(n61524), .ZN(n29410) );
  INV_X1 U33881 ( .A(n29410), .ZN(p_wishbone_bd_ram_n23223) );
  INV_X1 U33882 ( .A(n61523), .ZN(n29412) );
  INV_X1 U33883 ( .A(n29412), .ZN(p_wishbone_bd_ram_n23222) );
  INV_X1 U33884 ( .A(n61522), .ZN(n29414) );
  INV_X1 U33885 ( .A(n29414), .ZN(p_wishbone_bd_ram_n23221) );
  INV_X1 U33886 ( .A(n61521), .ZN(n29416) );
  INV_X1 U33887 ( .A(n29416), .ZN(p_wishbone_bd_ram_n23220) );
  INV_X1 U33888 ( .A(n61520), .ZN(n29418) );
  INV_X1 U33889 ( .A(n29418), .ZN(p_wishbone_bd_ram_n23219) );
  INV_X1 U33890 ( .A(n61519), .ZN(n29420) );
  INV_X1 U33891 ( .A(n29420), .ZN(p_wishbone_bd_ram_n23218) );
  INV_X1 U33892 ( .A(n61518), .ZN(n29422) );
  INV_X1 U33893 ( .A(n29422), .ZN(p_wishbone_bd_ram_n23217) );
  INV_X1 U33894 ( .A(n61517), .ZN(n29424) );
  INV_X1 U33895 ( .A(n29424), .ZN(p_wishbone_bd_ram_n23215) );
  INV_X1 U33896 ( .A(n61516), .ZN(n29426) );
  INV_X1 U33897 ( .A(n29426), .ZN(p_wishbone_bd_ram_n23213) );
  INV_X1 U33898 ( .A(n61515), .ZN(n29428) );
  INV_X1 U33899 ( .A(n29428), .ZN(p_wishbone_bd_ram_n23212) );
  INV_X1 U33900 ( .A(n61514), .ZN(n29430) );
  INV_X1 U33901 ( .A(n29430), .ZN(p_wishbone_bd_ram_n23210) );
  INV_X1 U33902 ( .A(n61513), .ZN(n29432) );
  INV_X1 U33903 ( .A(n29432), .ZN(p_wishbone_bd_ram_n23208) );
  INV_X1 U33904 ( .A(n61512), .ZN(n29434) );
  INV_X1 U33905 ( .A(n29434), .ZN(p_wishbone_bd_ram_n23207) );
  INV_X1 U33906 ( .A(n61511), .ZN(n29436) );
  INV_X1 U33907 ( .A(n29436), .ZN(p_wishbone_bd_ram_n23206) );
  INV_X1 U33908 ( .A(n61510), .ZN(n29438) );
  INV_X1 U33909 ( .A(n29438), .ZN(p_wishbone_bd_ram_n23205) );
  INV_X1 U33910 ( .A(n61509), .ZN(n29440) );
  INV_X1 U33911 ( .A(n29440), .ZN(p_wishbone_bd_ram_n23204) );
  INV_X1 U33912 ( .A(n61508), .ZN(n29442) );
  INV_X1 U33913 ( .A(n29442), .ZN(p_wishbone_bd_ram_n23203) );
  INV_X1 U33914 ( .A(n61507), .ZN(n29444) );
  INV_X1 U33915 ( .A(n29444), .ZN(p_wishbone_bd_ram_n23202) );
  INV_X1 U33916 ( .A(n61506), .ZN(n29446) );
  INV_X1 U33917 ( .A(n29446), .ZN(p_wishbone_bd_ram_n23201) );
  INV_X1 U33918 ( .A(n61505), .ZN(n29448) );
  INV_X1 U33919 ( .A(n29448), .ZN(p_wishbone_bd_ram_n23200) );
  INV_X1 U33920 ( .A(n61504), .ZN(n29450) );
  INV_X1 U33921 ( .A(n29450), .ZN(p_wishbone_bd_ram_n23199) );
  INV_X1 U33922 ( .A(n61503), .ZN(n29452) );
  INV_X1 U33923 ( .A(n29452), .ZN(p_wishbone_bd_ram_n23198) );
  INV_X1 U33924 ( .A(n61502), .ZN(n29454) );
  INV_X1 U33925 ( .A(n29454), .ZN(p_wishbone_bd_ram_n23197) );
  INV_X1 U33926 ( .A(n61501), .ZN(n29456) );
  INV_X1 U33927 ( .A(n29456), .ZN(p_wishbone_bd_ram_n23196) );
  INV_X1 U33928 ( .A(n61500), .ZN(n29458) );
  INV_X1 U33929 ( .A(n29458), .ZN(p_wishbone_bd_ram_n23195) );
  INV_X1 U33930 ( .A(n61499), .ZN(n29460) );
  INV_X1 U33931 ( .A(n29460), .ZN(p_wishbone_bd_ram_n23194) );
  INV_X1 U33932 ( .A(n61498), .ZN(n29462) );
  INV_X1 U33933 ( .A(n29462), .ZN(p_wishbone_bd_ram_n23193) );
  INV_X1 U33934 ( .A(n61497), .ZN(n29464) );
  INV_X1 U33935 ( .A(n29464), .ZN(p_wishbone_bd_ram_n23192) );
  INV_X1 U33936 ( .A(n61496), .ZN(n29466) );
  INV_X1 U33937 ( .A(n29466), .ZN(p_wishbone_bd_ram_n23191) );
  INV_X1 U33938 ( .A(n61495), .ZN(n29468) );
  INV_X1 U33939 ( .A(n29468), .ZN(p_wishbone_bd_ram_n23190) );
  INV_X1 U33940 ( .A(n61494), .ZN(n29470) );
  INV_X1 U33941 ( .A(n29470), .ZN(p_wishbone_bd_ram_n23189) );
  INV_X1 U33942 ( .A(n61493), .ZN(n29472) );
  INV_X1 U33943 ( .A(n29472), .ZN(p_wishbone_bd_ram_n23188) );
  INV_X1 U33944 ( .A(n61492), .ZN(n29474) );
  INV_X1 U33945 ( .A(n29474), .ZN(p_wishbone_bd_ram_n23187) );
  INV_X1 U33946 ( .A(n61491), .ZN(n29476) );
  INV_X1 U33947 ( .A(n29476), .ZN(p_wishbone_bd_ram_n23186) );
  INV_X1 U33948 ( .A(n61490), .ZN(n29478) );
  INV_X1 U33949 ( .A(n29478), .ZN(p_wishbone_bd_ram_n23185) );
  INV_X1 U33950 ( .A(n61489), .ZN(n29480) );
  INV_X1 U33951 ( .A(n29480), .ZN(p_wishbone_bd_ram_n23184) );
  INV_X1 U33952 ( .A(n61488), .ZN(n29482) );
  INV_X1 U33953 ( .A(n29482), .ZN(p_wishbone_bd_ram_n23183) );
  INV_X1 U33954 ( .A(n61487), .ZN(n29484) );
  INV_X1 U33955 ( .A(n29484), .ZN(p_wishbone_bd_ram_n23182) );
  INV_X1 U33956 ( .A(n61486), .ZN(n29486) );
  INV_X1 U33957 ( .A(n29486), .ZN(p_wishbone_bd_ram_n23181) );
  INV_X1 U33958 ( .A(n61485), .ZN(n29488) );
  INV_X1 U33959 ( .A(n29488), .ZN(p_wishbone_bd_ram_n23180) );
  INV_X1 U33960 ( .A(n61484), .ZN(n29490) );
  INV_X1 U33961 ( .A(n29490), .ZN(p_wishbone_bd_ram_n23179) );
  INV_X1 U33962 ( .A(n61483), .ZN(n29492) );
  INV_X1 U33963 ( .A(n29492), .ZN(p_wishbone_bd_ram_n23178) );
  INV_X1 U33964 ( .A(n61482), .ZN(n29494) );
  INV_X1 U33965 ( .A(n29494), .ZN(p_wishbone_bd_ram_n23177) );
  INV_X1 U33966 ( .A(n61481), .ZN(n29496) );
  INV_X1 U33967 ( .A(n29496), .ZN(p_wishbone_bd_ram_n23176) );
  INV_X1 U33968 ( .A(n61480), .ZN(n29498) );
  INV_X1 U33969 ( .A(n29498), .ZN(p_wishbone_bd_ram_n23175) );
  INV_X1 U33970 ( .A(n61479), .ZN(n29500) );
  INV_X1 U33971 ( .A(n29500), .ZN(p_wishbone_bd_ram_n23174) );
  INV_X1 U33972 ( .A(n61478), .ZN(n29502) );
  INV_X1 U33973 ( .A(n29502), .ZN(p_wishbone_bd_ram_n23173) );
  INV_X1 U33974 ( .A(n61477), .ZN(n29504) );
  INV_X1 U33975 ( .A(n29504), .ZN(p_wishbone_bd_ram_n23172) );
  INV_X1 U33976 ( .A(n61476), .ZN(n29506) );
  INV_X1 U33977 ( .A(n29506), .ZN(p_wishbone_bd_ram_n23171) );
  INV_X1 U33978 ( .A(n61475), .ZN(n29508) );
  INV_X1 U33979 ( .A(n29508), .ZN(p_wishbone_bd_ram_n23170) );
  INV_X1 U33980 ( .A(n61474), .ZN(n29510) );
  INV_X1 U33981 ( .A(n29510), .ZN(p_wishbone_bd_ram_n23169) );
  INV_X1 U33982 ( .A(n61473), .ZN(n29512) );
  INV_X1 U33983 ( .A(n29512), .ZN(p_wishbone_bd_ram_n23168) );
  INV_X1 U33984 ( .A(n61472), .ZN(n29514) );
  INV_X1 U33985 ( .A(n29514), .ZN(p_wishbone_bd_ram_n23167) );
  INV_X1 U33986 ( .A(n61471), .ZN(n29516) );
  INV_X1 U33987 ( .A(n29516), .ZN(p_wishbone_bd_ram_n23166) );
  INV_X1 U33988 ( .A(n61470), .ZN(n29518) );
  INV_X1 U33989 ( .A(n29518), .ZN(p_wishbone_bd_ram_n23165) );
  INV_X1 U33990 ( .A(n61469), .ZN(n29520) );
  INV_X1 U33991 ( .A(n29520), .ZN(p_wishbone_bd_ram_n23164) );
  INV_X1 U33992 ( .A(n61468), .ZN(n29522) );
  INV_X1 U33993 ( .A(n29522), .ZN(p_wishbone_bd_ram_n23163) );
  INV_X1 U33994 ( .A(n61467), .ZN(n29524) );
  INV_X1 U33995 ( .A(n29524), .ZN(p_wishbone_bd_ram_n23162) );
  INV_X1 U33996 ( .A(n61466), .ZN(n29526) );
  INV_X1 U33997 ( .A(n29526), .ZN(p_wishbone_bd_ram_n23161) );
  INV_X1 U33998 ( .A(n61465), .ZN(n29528) );
  INV_X1 U33999 ( .A(n29528), .ZN(p_wishbone_bd_ram_n23159) );
  INV_X1 U34000 ( .A(n61464), .ZN(n29530) );
  INV_X1 U34001 ( .A(n29530), .ZN(p_wishbone_bd_ram_n23157) );
  INV_X1 U34002 ( .A(n61463), .ZN(n29532) );
  INV_X1 U34003 ( .A(n29532), .ZN(p_wishbone_bd_ram_n23156) );
  INV_X1 U34004 ( .A(n61462), .ZN(n29534) );
  INV_X1 U34005 ( .A(n29534), .ZN(p_wishbone_bd_ram_n23154) );
  INV_X1 U34006 ( .A(n61461), .ZN(n29536) );
  INV_X1 U34007 ( .A(n29536), .ZN(p_wishbone_bd_ram_n23152) );
  INV_X1 U34008 ( .A(n61460), .ZN(n29538) );
  INV_X1 U34009 ( .A(n29538), .ZN(p_wishbone_bd_ram_n23151) );
  INV_X1 U34010 ( .A(n61459), .ZN(n29540) );
  INV_X1 U34011 ( .A(n29540), .ZN(p_wishbone_bd_ram_n23150) );
  INV_X1 U34012 ( .A(n61458), .ZN(n29542) );
  INV_X1 U34013 ( .A(n29542), .ZN(p_wishbone_bd_ram_n23149) );
  INV_X1 U34014 ( .A(n61457), .ZN(n29544) );
  INV_X1 U34015 ( .A(n29544), .ZN(p_wishbone_bd_ram_n23148) );
  INV_X1 U34016 ( .A(n61456), .ZN(n29546) );
  INV_X1 U34017 ( .A(n29546), .ZN(p_wishbone_bd_ram_n23147) );
  INV_X1 U34018 ( .A(n61455), .ZN(n29548) );
  INV_X1 U34019 ( .A(n29548), .ZN(p_wishbone_bd_ram_n23146) );
  INV_X1 U34020 ( .A(n61454), .ZN(n29550) );
  INV_X1 U34021 ( .A(n29550), .ZN(p_wishbone_bd_ram_n23145) );
  INV_X1 U34022 ( .A(n61453), .ZN(n29552) );
  INV_X1 U34023 ( .A(n29552), .ZN(p_wishbone_bd_ram_n23144) );
  INV_X1 U34024 ( .A(n61452), .ZN(n29554) );
  INV_X1 U34025 ( .A(n29554), .ZN(p_wishbone_bd_ram_n23143) );
  INV_X1 U34026 ( .A(n61451), .ZN(n29556) );
  INV_X1 U34027 ( .A(n29556), .ZN(p_wishbone_bd_ram_n23142) );
  INV_X1 U34028 ( .A(n61450), .ZN(n29558) );
  INV_X1 U34029 ( .A(n29558), .ZN(p_wishbone_bd_ram_n23141) );
  INV_X1 U34030 ( .A(n61449), .ZN(n29560) );
  INV_X1 U34031 ( .A(n29560), .ZN(p_wishbone_bd_ram_n23140) );
  INV_X1 U34032 ( .A(n61448), .ZN(n29562) );
  INV_X1 U34033 ( .A(n29562), .ZN(p_wishbone_bd_ram_n23139) );
  INV_X1 U34034 ( .A(n61447), .ZN(n29564) );
  INV_X1 U34035 ( .A(n29564), .ZN(p_wishbone_bd_ram_n23138) );
  INV_X1 U34036 ( .A(n61446), .ZN(n29566) );
  INV_X1 U34037 ( .A(n29566), .ZN(p_wishbone_bd_ram_n23137) );
  INV_X1 U34038 ( .A(n61445), .ZN(n29568) );
  INV_X1 U34039 ( .A(n29568), .ZN(p_wishbone_bd_ram_n23136) );
  INV_X1 U34040 ( .A(n61444), .ZN(n29570) );
  INV_X1 U34041 ( .A(n29570), .ZN(p_wishbone_bd_ram_n23135) );
  INV_X1 U34042 ( .A(n61443), .ZN(n29572) );
  INV_X1 U34043 ( .A(n29572), .ZN(p_wishbone_bd_ram_n23134) );
  INV_X1 U34044 ( .A(n61442), .ZN(n29574) );
  INV_X1 U34045 ( .A(n29574), .ZN(p_wishbone_bd_ram_n23133) );
  INV_X1 U34046 ( .A(n61441), .ZN(n29576) );
  INV_X1 U34047 ( .A(n29576), .ZN(p_wishbone_bd_ram_n23132) );
  INV_X1 U34048 ( .A(n61440), .ZN(n29578) );
  INV_X1 U34049 ( .A(n29578), .ZN(p_wishbone_bd_ram_n23131) );
  INV_X1 U34050 ( .A(n61439), .ZN(n29580) );
  INV_X1 U34051 ( .A(n29580), .ZN(p_wishbone_bd_ram_n23130) );
  INV_X1 U34052 ( .A(n61438), .ZN(n29582) );
  INV_X1 U34053 ( .A(n29582), .ZN(p_wishbone_bd_ram_n23129) );
  INV_X1 U34054 ( .A(n61437), .ZN(n29584) );
  INV_X1 U34055 ( .A(n29584), .ZN(p_wishbone_bd_ram_n23128) );
  INV_X1 U34056 ( .A(n61436), .ZN(n29586) );
  INV_X1 U34057 ( .A(n29586), .ZN(p_wishbone_bd_ram_n23127) );
  INV_X1 U34058 ( .A(n61435), .ZN(n29588) );
  INV_X1 U34059 ( .A(n29588), .ZN(p_wishbone_bd_ram_n23126) );
  INV_X1 U34060 ( .A(n61434), .ZN(n29590) );
  INV_X1 U34061 ( .A(n29590), .ZN(p_wishbone_bd_ram_n23125) );
  INV_X1 U34062 ( .A(n61433), .ZN(n29592) );
  INV_X1 U34063 ( .A(n29592), .ZN(p_wishbone_bd_ram_n23124) );
  INV_X1 U34064 ( .A(n61432), .ZN(n29594) );
  INV_X1 U34065 ( .A(n29594), .ZN(p_wishbone_bd_ram_n23123) );
  INV_X1 U34066 ( .A(n61431), .ZN(n29596) );
  INV_X1 U34067 ( .A(n29596), .ZN(p_wishbone_bd_ram_n23122) );
  INV_X1 U34068 ( .A(n61430), .ZN(n29598) );
  INV_X1 U34069 ( .A(n29598), .ZN(p_wishbone_bd_ram_n23121) );
  INV_X1 U34070 ( .A(n61429), .ZN(n29600) );
  INV_X1 U34071 ( .A(n29600), .ZN(p_wishbone_bd_ram_n23120) );
  INV_X1 U34072 ( .A(n61428), .ZN(n29602) );
  INV_X1 U34073 ( .A(n29602), .ZN(p_wishbone_bd_ram_n23119) );
  INV_X1 U34074 ( .A(n61427), .ZN(n29604) );
  INV_X1 U34075 ( .A(n29604), .ZN(p_wishbone_bd_ram_n23118) );
  INV_X1 U34076 ( .A(n61426), .ZN(n29606) );
  INV_X1 U34077 ( .A(n29606), .ZN(p_wishbone_bd_ram_n23117) );
  INV_X1 U34078 ( .A(n61425), .ZN(n29608) );
  INV_X1 U34079 ( .A(n29608), .ZN(p_wishbone_bd_ram_n23116) );
  INV_X1 U34080 ( .A(n61424), .ZN(n29610) );
  INV_X1 U34081 ( .A(n29610), .ZN(p_wishbone_bd_ram_n23115) );
  INV_X1 U34082 ( .A(n61423), .ZN(n29612) );
  INV_X1 U34083 ( .A(n29612), .ZN(p_wishbone_bd_ram_n23114) );
  INV_X1 U34084 ( .A(n61422), .ZN(n29614) );
  INV_X1 U34085 ( .A(n29614), .ZN(p_wishbone_bd_ram_n23113) );
  INV_X1 U34086 ( .A(n61421), .ZN(n29616) );
  INV_X1 U34087 ( .A(n29616), .ZN(p_wishbone_bd_ram_n23112) );
  INV_X1 U34088 ( .A(n61420), .ZN(n29618) );
  INV_X1 U34089 ( .A(n29618), .ZN(p_wishbone_bd_ram_n23111) );
  INV_X1 U34090 ( .A(n61419), .ZN(n29620) );
  INV_X1 U34091 ( .A(n29620), .ZN(p_wishbone_bd_ram_n23110) );
  INV_X1 U34092 ( .A(n61418), .ZN(n29622) );
  INV_X1 U34093 ( .A(n29622), .ZN(p_wishbone_bd_ram_n23109) );
  INV_X1 U34094 ( .A(n61417), .ZN(n29624) );
  INV_X1 U34095 ( .A(n29624), .ZN(p_wishbone_bd_ram_n23108) );
  INV_X1 U34096 ( .A(n61416), .ZN(n29626) );
  INV_X1 U34097 ( .A(n29626), .ZN(p_wishbone_bd_ram_n23107) );
  INV_X1 U34098 ( .A(n61415), .ZN(n29628) );
  INV_X1 U34099 ( .A(n29628), .ZN(p_wishbone_bd_ram_n23106) );
  INV_X1 U34100 ( .A(n61414), .ZN(n29630) );
  INV_X1 U34101 ( .A(n29630), .ZN(p_wishbone_bd_ram_n23105) );
  INV_X1 U34102 ( .A(n61413), .ZN(n29632) );
  INV_X1 U34103 ( .A(n29632), .ZN(p_wishbone_bd_ram_n23104) );
  INV_X1 U34104 ( .A(n61412), .ZN(n29634) );
  INV_X1 U34105 ( .A(n29634), .ZN(p_wishbone_bd_ram_n23103) );
  INV_X1 U34106 ( .A(n61411), .ZN(n29636) );
  INV_X1 U34107 ( .A(n29636), .ZN(p_wishbone_bd_ram_n23102) );
  INV_X1 U34108 ( .A(n61410), .ZN(n29638) );
  INV_X1 U34109 ( .A(n29638), .ZN(p_wishbone_bd_ram_n23101) );
  INV_X1 U34110 ( .A(n61409), .ZN(n29640) );
  INV_X1 U34111 ( .A(n29640), .ZN(p_wishbone_bd_ram_n23100) );
  INV_X1 U34112 ( .A(n61408), .ZN(n29642) );
  INV_X1 U34113 ( .A(n29642), .ZN(p_wishbone_bd_ram_n23099) );
  INV_X1 U34114 ( .A(n61407), .ZN(n29644) );
  INV_X1 U34115 ( .A(n29644), .ZN(p_wishbone_bd_ram_n23098) );
  INV_X1 U34116 ( .A(n61406), .ZN(n29646) );
  INV_X1 U34117 ( .A(n29646), .ZN(p_wishbone_bd_ram_n23097) );
  INV_X1 U34118 ( .A(n61405), .ZN(n29648) );
  INV_X1 U34119 ( .A(n29648), .ZN(p_wishbone_bd_ram_n23096) );
  INV_X1 U34120 ( .A(n61404), .ZN(n29650) );
  INV_X1 U34121 ( .A(n29650), .ZN(p_wishbone_bd_ram_n23095) );
  INV_X1 U34122 ( .A(n61403), .ZN(n29652) );
  INV_X1 U34123 ( .A(n29652), .ZN(p_wishbone_bd_ram_n23094) );
  INV_X1 U34124 ( .A(n61402), .ZN(n29654) );
  INV_X1 U34125 ( .A(n29654), .ZN(p_wishbone_bd_ram_n23093) );
  INV_X1 U34126 ( .A(n61401), .ZN(n29656) );
  INV_X1 U34127 ( .A(n29656), .ZN(p_wishbone_bd_ram_n23092) );
  INV_X1 U34128 ( .A(n61400), .ZN(n29658) );
  INV_X1 U34129 ( .A(n29658), .ZN(p_wishbone_bd_ram_n23091) );
  INV_X1 U34130 ( .A(n61399), .ZN(n29660) );
  INV_X1 U34131 ( .A(n29660), .ZN(p_wishbone_bd_ram_n23090) );
  INV_X1 U34132 ( .A(n61398), .ZN(n29662) );
  INV_X1 U34133 ( .A(n29662), .ZN(p_wishbone_bd_ram_n23089) );
  INV_X1 U34134 ( .A(n61397), .ZN(n29664) );
  INV_X1 U34135 ( .A(n29664), .ZN(p_wishbone_bd_ram_n23087) );
  INV_X1 U34136 ( .A(n61396), .ZN(n29666) );
  INV_X1 U34137 ( .A(n29666), .ZN(p_wishbone_bd_ram_n23085) );
  INV_X1 U34138 ( .A(n61395), .ZN(n29668) );
  INV_X1 U34139 ( .A(n29668), .ZN(p_wishbone_bd_ram_n23084) );
  INV_X1 U34140 ( .A(n61394), .ZN(n29670) );
  INV_X1 U34141 ( .A(n29670), .ZN(p_wishbone_bd_ram_n23082) );
  INV_X1 U34142 ( .A(n61393), .ZN(n29672) );
  INV_X1 U34143 ( .A(n29672), .ZN(p_wishbone_bd_ram_n23080) );
  INV_X1 U34144 ( .A(n61392), .ZN(n29674) );
  INV_X1 U34145 ( .A(n29674), .ZN(p_wishbone_bd_ram_n23079) );
  INV_X1 U34146 ( .A(n61391), .ZN(n29676) );
  INV_X1 U34147 ( .A(n29676), .ZN(p_wishbone_bd_ram_n23078) );
  INV_X1 U34148 ( .A(n61390), .ZN(n29678) );
  INV_X1 U34149 ( .A(n29678), .ZN(p_wishbone_bd_ram_n23077) );
  INV_X1 U34150 ( .A(n61389), .ZN(n29680) );
  INV_X1 U34151 ( .A(n29680), .ZN(p_wishbone_bd_ram_n23076) );
  INV_X1 U34152 ( .A(n61388), .ZN(n29682) );
  INV_X1 U34153 ( .A(n29682), .ZN(p_wishbone_bd_ram_n23075) );
  INV_X1 U34154 ( .A(n61387), .ZN(n29684) );
  INV_X1 U34155 ( .A(n29684), .ZN(p_wishbone_bd_ram_n23074) );
  INV_X1 U34156 ( .A(n61386), .ZN(n29686) );
  INV_X1 U34157 ( .A(n29686), .ZN(p_wishbone_bd_ram_n23073) );
  INV_X1 U34158 ( .A(n61385), .ZN(n29688) );
  INV_X1 U34159 ( .A(n29688), .ZN(p_wishbone_bd_ram_n23072) );
  INV_X1 U34160 ( .A(n61384), .ZN(n29690) );
  INV_X1 U34161 ( .A(n29690), .ZN(p_wishbone_bd_ram_n23071) );
  INV_X1 U34162 ( .A(n61383), .ZN(n29692) );
  INV_X1 U34163 ( .A(n29692), .ZN(p_wishbone_bd_ram_n23070) );
  INV_X1 U34164 ( .A(n61382), .ZN(n29694) );
  INV_X1 U34165 ( .A(n29694), .ZN(p_wishbone_bd_ram_n23069) );
  INV_X1 U34166 ( .A(n61381), .ZN(n29696) );
  INV_X1 U34167 ( .A(n29696), .ZN(p_wishbone_bd_ram_n23068) );
  INV_X1 U34168 ( .A(n61380), .ZN(n29698) );
  INV_X1 U34169 ( .A(n29698), .ZN(p_wishbone_bd_ram_n23067) );
  INV_X1 U34170 ( .A(n61379), .ZN(n29700) );
  INV_X1 U34171 ( .A(n29700), .ZN(p_wishbone_bd_ram_n23066) );
  INV_X1 U34172 ( .A(n61378), .ZN(n29702) );
  INV_X1 U34173 ( .A(n29702), .ZN(p_wishbone_bd_ram_n23065) );
  INV_X1 U34174 ( .A(n61377), .ZN(n29704) );
  INV_X1 U34175 ( .A(n29704), .ZN(p_wishbone_bd_ram_n23064) );
  INV_X1 U34176 ( .A(n61376), .ZN(n29706) );
  INV_X1 U34177 ( .A(n29706), .ZN(p_wishbone_bd_ram_n23063) );
  INV_X1 U34178 ( .A(n61375), .ZN(n29708) );
  INV_X1 U34179 ( .A(n29708), .ZN(p_wishbone_bd_ram_n23062) );
  INV_X1 U34180 ( .A(n61374), .ZN(n29710) );
  INV_X1 U34181 ( .A(n29710), .ZN(p_wishbone_bd_ram_n23061) );
  INV_X1 U34182 ( .A(n61373), .ZN(n29712) );
  INV_X1 U34183 ( .A(n29712), .ZN(p_wishbone_bd_ram_n23060) );
  INV_X1 U34184 ( .A(n61372), .ZN(n29714) );
  INV_X1 U34185 ( .A(n29714), .ZN(p_wishbone_bd_ram_n23059) );
  INV_X1 U34186 ( .A(n61371), .ZN(n29716) );
  INV_X1 U34187 ( .A(n29716), .ZN(p_wishbone_bd_ram_n23058) );
  INV_X1 U34188 ( .A(n61370), .ZN(n29718) );
  INV_X1 U34189 ( .A(n29718), .ZN(p_wishbone_bd_ram_n23057) );
  INV_X1 U34190 ( .A(n61369), .ZN(n29720) );
  INV_X1 U34191 ( .A(n29720), .ZN(p_wishbone_bd_ram_n23056) );
  INV_X1 U34192 ( .A(n61368), .ZN(n29722) );
  INV_X1 U34193 ( .A(n29722), .ZN(p_wishbone_bd_ram_n23055) );
  INV_X1 U34194 ( .A(n61367), .ZN(n29724) );
  INV_X1 U34195 ( .A(n29724), .ZN(p_wishbone_bd_ram_n23054) );
  INV_X1 U34196 ( .A(n61366), .ZN(n29726) );
  INV_X1 U34197 ( .A(n29726), .ZN(p_wishbone_bd_ram_n23053) );
  INV_X1 U34198 ( .A(n61365), .ZN(n29728) );
  INV_X1 U34199 ( .A(n29728), .ZN(p_wishbone_bd_ram_n23052) );
  INV_X1 U34200 ( .A(n61364), .ZN(n29730) );
  INV_X1 U34201 ( .A(n29730), .ZN(p_wishbone_bd_ram_n23051) );
  INV_X1 U34202 ( .A(n61363), .ZN(n29732) );
  INV_X1 U34203 ( .A(n29732), .ZN(p_wishbone_bd_ram_n23050) );
  INV_X1 U34204 ( .A(n61362), .ZN(n29734) );
  INV_X1 U34205 ( .A(n29734), .ZN(p_wishbone_bd_ram_n23049) );
  INV_X1 U34206 ( .A(n61361), .ZN(n29736) );
  INV_X1 U34207 ( .A(n29736), .ZN(p_wishbone_bd_ram_n23048) );
  INV_X1 U34208 ( .A(n61360), .ZN(n29738) );
  INV_X1 U34209 ( .A(n29738), .ZN(p_wishbone_bd_ram_n23047) );
  INV_X1 U34210 ( .A(n61359), .ZN(n29740) );
  INV_X1 U34211 ( .A(n29740), .ZN(p_wishbone_bd_ram_n23046) );
  INV_X1 U34212 ( .A(n61358), .ZN(n29742) );
  INV_X1 U34213 ( .A(n29742), .ZN(p_wishbone_bd_ram_n23045) );
  INV_X1 U34214 ( .A(n61357), .ZN(n29744) );
  INV_X1 U34215 ( .A(n29744), .ZN(p_wishbone_bd_ram_n23044) );
  INV_X1 U34216 ( .A(n61356), .ZN(n29746) );
  INV_X1 U34217 ( .A(n29746), .ZN(p_wishbone_bd_ram_n23043) );
  INV_X1 U34218 ( .A(n61355), .ZN(n29748) );
  INV_X1 U34219 ( .A(n29748), .ZN(p_wishbone_bd_ram_n23042) );
  INV_X1 U34220 ( .A(n61354), .ZN(n29750) );
  INV_X1 U34221 ( .A(n29750), .ZN(p_wishbone_bd_ram_n23041) );
  INV_X1 U34222 ( .A(n61353), .ZN(n29752) );
  INV_X1 U34223 ( .A(n29752), .ZN(p_wishbone_bd_ram_n23040) );
  INV_X1 U34224 ( .A(n61352), .ZN(n29754) );
  INV_X1 U34225 ( .A(n29754), .ZN(p_wishbone_bd_ram_n23039) );
  INV_X1 U34226 ( .A(n61351), .ZN(n29756) );
  INV_X1 U34227 ( .A(n29756), .ZN(p_wishbone_bd_ram_n23038) );
  INV_X1 U34228 ( .A(n61350), .ZN(n29758) );
  INV_X1 U34229 ( .A(n29758), .ZN(p_wishbone_bd_ram_n23037) );
  INV_X1 U34230 ( .A(n61349), .ZN(n29760) );
  INV_X1 U34231 ( .A(n29760), .ZN(p_wishbone_bd_ram_n23036) );
  INV_X1 U34232 ( .A(n61348), .ZN(n29762) );
  INV_X1 U34233 ( .A(n29762), .ZN(p_wishbone_bd_ram_n23035) );
  INV_X1 U34234 ( .A(n61347), .ZN(n29764) );
  INV_X1 U34235 ( .A(n29764), .ZN(p_wishbone_bd_ram_n23034) );
  INV_X1 U34236 ( .A(n61346), .ZN(n29766) );
  INV_X1 U34237 ( .A(n29766), .ZN(p_wishbone_bd_ram_n23033) );
  INV_X1 U34238 ( .A(n61345), .ZN(n29768) );
  INV_X1 U34239 ( .A(n29768), .ZN(p_wishbone_bd_ram_n23032) );
  INV_X1 U34240 ( .A(n61344), .ZN(n29770) );
  INV_X1 U34241 ( .A(n29770), .ZN(p_wishbone_bd_ram_n23031) );
  INV_X1 U34242 ( .A(n61343), .ZN(n29772) );
  INV_X1 U34243 ( .A(n29772), .ZN(p_wishbone_bd_ram_n23030) );
  INV_X1 U34244 ( .A(n61342), .ZN(n29774) );
  INV_X1 U34245 ( .A(n29774), .ZN(p_wishbone_bd_ram_n23029) );
  INV_X1 U34246 ( .A(n61341), .ZN(n29776) );
  INV_X1 U34247 ( .A(n29776), .ZN(p_wishbone_bd_ram_n23028) );
  INV_X1 U34248 ( .A(n61340), .ZN(n29778) );
  INV_X1 U34249 ( .A(n29778), .ZN(p_wishbone_bd_ram_n23027) );
  INV_X1 U34250 ( .A(n61339), .ZN(n29780) );
  INV_X1 U34251 ( .A(n29780), .ZN(p_wishbone_bd_ram_n23026) );
  INV_X1 U34252 ( .A(n61338), .ZN(n29782) );
  INV_X1 U34253 ( .A(n29782), .ZN(p_wishbone_bd_ram_n23025) );
  INV_X1 U34254 ( .A(n61337), .ZN(n29784) );
  INV_X1 U34255 ( .A(n29784), .ZN(p_wishbone_bd_ram_n23023) );
  INV_X1 U34256 ( .A(n61336), .ZN(n29786) );
  INV_X1 U34257 ( .A(n29786), .ZN(p_wishbone_bd_ram_n23021) );
  INV_X1 U34258 ( .A(n61335), .ZN(n29788) );
  INV_X1 U34259 ( .A(n29788), .ZN(p_wishbone_bd_ram_n23020) );
  INV_X1 U34260 ( .A(n61334), .ZN(n29790) );
  INV_X1 U34261 ( .A(n29790), .ZN(p_wishbone_bd_ram_n23018) );
  INV_X1 U34262 ( .A(n61333), .ZN(n29792) );
  INV_X1 U34263 ( .A(n29792), .ZN(p_wishbone_bd_ram_n23016) );
  INV_X1 U34264 ( .A(n61332), .ZN(n29794) );
  INV_X1 U34265 ( .A(n29794), .ZN(p_wishbone_bd_ram_n23015) );
  INV_X1 U34266 ( .A(n61331), .ZN(n29796) );
  INV_X1 U34267 ( .A(n29796), .ZN(p_wishbone_bd_ram_n23014) );
  INV_X1 U34268 ( .A(n61330), .ZN(n29798) );
  INV_X1 U34269 ( .A(n29798), .ZN(p_wishbone_bd_ram_n23013) );
  INV_X1 U34270 ( .A(n61329), .ZN(n29800) );
  INV_X1 U34271 ( .A(n29800), .ZN(p_wishbone_bd_ram_n23012) );
  INV_X1 U34272 ( .A(n61328), .ZN(n29802) );
  INV_X1 U34273 ( .A(n29802), .ZN(p_wishbone_bd_ram_n23011) );
  INV_X1 U34274 ( .A(n61327), .ZN(n29804) );
  INV_X1 U34275 ( .A(n29804), .ZN(p_wishbone_bd_ram_n23010) );
  INV_X1 U34276 ( .A(n61326), .ZN(n29806) );
  INV_X1 U34277 ( .A(n29806), .ZN(p_wishbone_bd_ram_n23009) );
  INV_X1 U34278 ( .A(n61325), .ZN(n29808) );
  INV_X1 U34279 ( .A(n29808), .ZN(p_wishbone_bd_ram_n23008) );
  INV_X1 U34280 ( .A(n61324), .ZN(n29810) );
  INV_X1 U34281 ( .A(n29810), .ZN(p_wishbone_bd_ram_n23007) );
  INV_X1 U34282 ( .A(n61323), .ZN(n29812) );
  INV_X1 U34283 ( .A(n29812), .ZN(p_wishbone_bd_ram_n23006) );
  INV_X1 U34284 ( .A(n61322), .ZN(n29814) );
  INV_X1 U34285 ( .A(n29814), .ZN(p_wishbone_bd_ram_n23005) );
  INV_X1 U34286 ( .A(n61321), .ZN(n29816) );
  INV_X1 U34287 ( .A(n29816), .ZN(p_wishbone_bd_ram_n23004) );
  INV_X1 U34288 ( .A(n61320), .ZN(n29818) );
  INV_X1 U34289 ( .A(n29818), .ZN(p_wishbone_bd_ram_n23003) );
  INV_X1 U34290 ( .A(n61319), .ZN(n29820) );
  INV_X1 U34291 ( .A(n29820), .ZN(p_wishbone_bd_ram_n23002) );
  INV_X1 U34292 ( .A(n61318), .ZN(n29822) );
  INV_X1 U34293 ( .A(n29822), .ZN(p_wishbone_bd_ram_n23001) );
  INV_X1 U34294 ( .A(n61317), .ZN(n29824) );
  INV_X1 U34295 ( .A(n29824), .ZN(p_wishbone_bd_ram_n23000) );
  INV_X1 U34296 ( .A(n61316), .ZN(n29826) );
  INV_X1 U34297 ( .A(n29826), .ZN(p_wishbone_bd_ram_n22999) );
  INV_X1 U34298 ( .A(n61315), .ZN(n29828) );
  INV_X1 U34299 ( .A(n29828), .ZN(p_wishbone_bd_ram_n22998) );
  INV_X1 U34300 ( .A(n61314), .ZN(n29830) );
  INV_X1 U34301 ( .A(n29830), .ZN(p_wishbone_bd_ram_n22997) );
  INV_X1 U34302 ( .A(n61313), .ZN(n29832) );
  INV_X1 U34303 ( .A(n29832), .ZN(p_wishbone_bd_ram_n22996) );
  INV_X1 U34304 ( .A(n61312), .ZN(n29834) );
  INV_X1 U34305 ( .A(n29834), .ZN(p_wishbone_bd_ram_n22995) );
  INV_X1 U34306 ( .A(n61311), .ZN(n29836) );
  INV_X1 U34307 ( .A(n29836), .ZN(p_wishbone_bd_ram_n22994) );
  INV_X1 U34308 ( .A(n61310), .ZN(n29838) );
  INV_X1 U34309 ( .A(n29838), .ZN(p_wishbone_bd_ram_n22993) );
  INV_X1 U34310 ( .A(n61309), .ZN(n29840) );
  INV_X1 U34311 ( .A(n29840), .ZN(p_wishbone_bd_ram_n22992) );
  INV_X1 U34312 ( .A(n61308), .ZN(n29842) );
  INV_X1 U34313 ( .A(n29842), .ZN(p_wishbone_bd_ram_n22991) );
  INV_X1 U34314 ( .A(n61307), .ZN(n29844) );
  INV_X1 U34315 ( .A(n29844), .ZN(p_wishbone_bd_ram_n22990) );
  INV_X1 U34316 ( .A(n61306), .ZN(n29846) );
  INV_X1 U34317 ( .A(n29846), .ZN(p_wishbone_bd_ram_n22989) );
  INV_X1 U34318 ( .A(n61305), .ZN(n29848) );
  INV_X1 U34319 ( .A(n29848), .ZN(p_wishbone_bd_ram_n22988) );
  INV_X1 U34320 ( .A(n61304), .ZN(n29850) );
  INV_X1 U34321 ( .A(n29850), .ZN(p_wishbone_bd_ram_n22987) );
  INV_X1 U34322 ( .A(n61303), .ZN(n29852) );
  INV_X1 U34323 ( .A(n29852), .ZN(p_wishbone_bd_ram_n22986) );
  INV_X1 U34324 ( .A(n61302), .ZN(n29854) );
  INV_X1 U34325 ( .A(n29854), .ZN(p_wishbone_bd_ram_n22985) );
  INV_X1 U34326 ( .A(n61301), .ZN(n29856) );
  INV_X1 U34327 ( .A(n29856), .ZN(p_wishbone_bd_ram_n22984) );
  INV_X1 U34328 ( .A(n61300), .ZN(n29858) );
  INV_X1 U34329 ( .A(n29858), .ZN(p_wishbone_bd_ram_n22983) );
  INV_X1 U34330 ( .A(n61299), .ZN(n29860) );
  INV_X1 U34331 ( .A(n29860), .ZN(p_wishbone_bd_ram_n22982) );
  INV_X1 U34332 ( .A(n61298), .ZN(n29862) );
  INV_X1 U34333 ( .A(n29862), .ZN(p_wishbone_bd_ram_n22981) );
  INV_X1 U34334 ( .A(n61297), .ZN(n29864) );
  INV_X1 U34335 ( .A(n29864), .ZN(p_wishbone_bd_ram_n22980) );
  INV_X1 U34336 ( .A(n61296), .ZN(n29866) );
  INV_X1 U34337 ( .A(n29866), .ZN(p_wishbone_bd_ram_n22979) );
  INV_X1 U34338 ( .A(n61295), .ZN(n29868) );
  INV_X1 U34339 ( .A(n29868), .ZN(p_wishbone_bd_ram_n22978) );
  INV_X1 U34340 ( .A(n61294), .ZN(n29870) );
  INV_X1 U34341 ( .A(n29870), .ZN(p_wishbone_bd_ram_n22977) );
  INV_X1 U34342 ( .A(n61293), .ZN(n29872) );
  INV_X1 U34343 ( .A(n29872), .ZN(p_wishbone_bd_ram_n22975) );
  INV_X1 U34344 ( .A(n61292), .ZN(n29874) );
  INV_X1 U34345 ( .A(n29874), .ZN(p_wishbone_bd_ram_n22973) );
  INV_X1 U34346 ( .A(n61291), .ZN(n29876) );
  INV_X1 U34347 ( .A(n29876), .ZN(p_wishbone_bd_ram_n22972) );
  INV_X1 U34348 ( .A(n61290), .ZN(n29878) );
  INV_X1 U34349 ( .A(n29878), .ZN(p_wishbone_bd_ram_n22970) );
  INV_X1 U34350 ( .A(n61289), .ZN(n29880) );
  INV_X1 U34351 ( .A(n29880), .ZN(p_wishbone_bd_ram_n22968) );
  INV_X1 U34352 ( .A(n61288), .ZN(n29882) );
  INV_X1 U34353 ( .A(n29882), .ZN(p_wishbone_bd_ram_n22967) );
  INV_X1 U34354 ( .A(n61287), .ZN(n29884) );
  INV_X1 U34355 ( .A(n29884), .ZN(p_wishbone_bd_ram_n22966) );
  INV_X1 U34356 ( .A(n61286), .ZN(n29886) );
  INV_X1 U34357 ( .A(n29886), .ZN(p_wishbone_bd_ram_n22965) );
  INV_X1 U34358 ( .A(n61285), .ZN(n29888) );
  INV_X1 U34359 ( .A(n29888), .ZN(p_wishbone_bd_ram_n22964) );
  INV_X1 U34360 ( .A(n61284), .ZN(n29890) );
  INV_X1 U34361 ( .A(n29890), .ZN(p_wishbone_bd_ram_n22963) );
  INV_X1 U34362 ( .A(n61283), .ZN(n29892) );
  INV_X1 U34363 ( .A(n29892), .ZN(p_wishbone_bd_ram_n22962) );
  INV_X1 U34364 ( .A(n61282), .ZN(n29894) );
  INV_X1 U34365 ( .A(n29894), .ZN(p_wishbone_bd_ram_n22961) );
  INV_X1 U34366 ( .A(n61281), .ZN(n29896) );
  INV_X1 U34367 ( .A(n29896), .ZN(p_wishbone_bd_ram_n22960) );
  INV_X1 U34368 ( .A(n61280), .ZN(n29898) );
  INV_X1 U34369 ( .A(n29898), .ZN(p_wishbone_bd_ram_n22959) );
  INV_X1 U34370 ( .A(n61279), .ZN(n29900) );
  INV_X1 U34371 ( .A(n29900), .ZN(p_wishbone_bd_ram_n22958) );
  INV_X1 U34372 ( .A(n61278), .ZN(n29902) );
  INV_X1 U34373 ( .A(n29902), .ZN(p_wishbone_bd_ram_n22957) );
  INV_X1 U34374 ( .A(n61277), .ZN(n29904) );
  INV_X1 U34375 ( .A(n29904), .ZN(p_wishbone_bd_ram_n22956) );
  INV_X1 U34376 ( .A(n61276), .ZN(n29906) );
  INV_X1 U34377 ( .A(n29906), .ZN(p_wishbone_bd_ram_n22955) );
  INV_X1 U34378 ( .A(n61275), .ZN(n29908) );
  INV_X1 U34379 ( .A(n29908), .ZN(p_wishbone_bd_ram_n22954) );
  INV_X1 U34380 ( .A(n61274), .ZN(n29910) );
  INV_X1 U34381 ( .A(n29910), .ZN(p_wishbone_bd_ram_n22953) );
  INV_X1 U34382 ( .A(n61273), .ZN(n29912) );
  INV_X1 U34383 ( .A(n29912), .ZN(p_wishbone_bd_ram_n22951) );
  INV_X1 U34384 ( .A(n61272), .ZN(n29914) );
  INV_X1 U34385 ( .A(n29914), .ZN(p_wishbone_bd_ram_n22949) );
  INV_X1 U34386 ( .A(n61271), .ZN(n29916) );
  INV_X1 U34387 ( .A(n29916), .ZN(p_wishbone_bd_ram_n22948) );
  INV_X1 U34388 ( .A(n61270), .ZN(n29918) );
  INV_X1 U34389 ( .A(n29918), .ZN(p_wishbone_bd_ram_n22946) );
  INV_X1 U34390 ( .A(n61269), .ZN(n29920) );
  INV_X1 U34391 ( .A(n29920), .ZN(p_wishbone_bd_ram_n22944) );
  INV_X1 U34392 ( .A(n61268), .ZN(n29922) );
  INV_X1 U34393 ( .A(n29922), .ZN(p_wishbone_bd_ram_n22943) );
  INV_X1 U34394 ( .A(n61267), .ZN(n29924) );
  INV_X1 U34395 ( .A(n29924), .ZN(p_wishbone_bd_ram_n22942) );
  INV_X1 U34396 ( .A(n61266), .ZN(n29926) );
  INV_X1 U34397 ( .A(n29926), .ZN(p_wishbone_bd_ram_n22941) );
  INV_X1 U34398 ( .A(n61265), .ZN(n29928) );
  INV_X1 U34399 ( .A(n29928), .ZN(p_wishbone_bd_ram_n22940) );
  INV_X1 U34400 ( .A(n61264), .ZN(n29930) );
  INV_X1 U34401 ( .A(n29930), .ZN(p_wishbone_bd_ram_n22939) );
  INV_X1 U34402 ( .A(n61263), .ZN(n29932) );
  INV_X1 U34403 ( .A(n29932), .ZN(p_wishbone_bd_ram_n22938) );
  INV_X1 U34404 ( .A(n61262), .ZN(n29934) );
  INV_X1 U34405 ( .A(n29934), .ZN(p_wishbone_bd_ram_n22937) );
  INV_X1 U34406 ( .A(n61261), .ZN(n29936) );
  INV_X1 U34407 ( .A(n29936), .ZN(p_wishbone_bd_ram_n22936) );
  INV_X1 U34408 ( .A(n61260), .ZN(n29938) );
  INV_X1 U34409 ( .A(n29938), .ZN(p_wishbone_bd_ram_n22935) );
  INV_X1 U34410 ( .A(n61259), .ZN(n29940) );
  INV_X1 U34411 ( .A(n29940), .ZN(p_wishbone_bd_ram_n22934) );
  INV_X1 U34412 ( .A(n61258), .ZN(n29942) );
  INV_X1 U34413 ( .A(n29942), .ZN(p_wishbone_bd_ram_n22933) );
  INV_X1 U34414 ( .A(n61257), .ZN(n29944) );
  INV_X1 U34415 ( .A(n29944), .ZN(p_wishbone_bd_ram_n22932) );
  INV_X1 U34416 ( .A(n61256), .ZN(n29946) );
  INV_X1 U34417 ( .A(n29946), .ZN(p_wishbone_bd_ram_n22931) );
  INV_X1 U34418 ( .A(n61255), .ZN(n29948) );
  INV_X1 U34419 ( .A(n29948), .ZN(p_wishbone_bd_ram_n22930) );
  INV_X1 U34420 ( .A(n61254), .ZN(n29950) );
  INV_X1 U34421 ( .A(n29950), .ZN(p_wishbone_bd_ram_n22929) );
  INV_X1 U34422 ( .A(n61253), .ZN(n29952) );
  INV_X1 U34423 ( .A(n29952), .ZN(p_wishbone_bd_ram_n22928) );
  INV_X1 U34424 ( .A(n61252), .ZN(n29954) );
  INV_X1 U34425 ( .A(n29954), .ZN(p_wishbone_bd_ram_n22927) );
  INV_X1 U34426 ( .A(n61251), .ZN(n29956) );
  INV_X1 U34427 ( .A(n29956), .ZN(p_wishbone_bd_ram_n22926) );
  INV_X1 U34428 ( .A(n61250), .ZN(n29958) );
  INV_X1 U34429 ( .A(n29958), .ZN(p_wishbone_bd_ram_n22925) );
  INV_X1 U34430 ( .A(n61249), .ZN(n29960) );
  INV_X1 U34431 ( .A(n29960), .ZN(p_wishbone_bd_ram_n22924) );
  INV_X1 U34432 ( .A(n61248), .ZN(n29962) );
  INV_X1 U34433 ( .A(n29962), .ZN(p_wishbone_bd_ram_n22923) );
  INV_X1 U34434 ( .A(n61247), .ZN(n29964) );
  INV_X1 U34435 ( .A(n29964), .ZN(p_wishbone_bd_ram_n22922) );
  INV_X1 U34436 ( .A(n61246), .ZN(n29966) );
  INV_X1 U34437 ( .A(n29966), .ZN(p_wishbone_bd_ram_n22921) );
  INV_X1 U34438 ( .A(n61245), .ZN(n29968) );
  INV_X1 U34439 ( .A(n29968), .ZN(p_wishbone_bd_ram_n22920) );
  INV_X1 U34440 ( .A(n61244), .ZN(n29970) );
  INV_X1 U34441 ( .A(n29970), .ZN(p_wishbone_bd_ram_n22919) );
  INV_X1 U34442 ( .A(n61243), .ZN(n29972) );
  INV_X1 U34443 ( .A(n29972), .ZN(p_wishbone_bd_ram_n22918) );
  INV_X1 U34444 ( .A(n61242), .ZN(n29974) );
  INV_X1 U34445 ( .A(n29974), .ZN(p_wishbone_bd_ram_n22917) );
  INV_X1 U34446 ( .A(n61241), .ZN(n29976) );
  INV_X1 U34447 ( .A(n29976), .ZN(p_wishbone_bd_ram_n22916) );
  INV_X1 U34448 ( .A(n61240), .ZN(n29978) );
  INV_X1 U34449 ( .A(n29978), .ZN(p_wishbone_bd_ram_n22915) );
  INV_X1 U34450 ( .A(n61239), .ZN(n29980) );
  INV_X1 U34451 ( .A(n29980), .ZN(p_wishbone_bd_ram_n22914) );
  INV_X1 U34452 ( .A(n61238), .ZN(n29982) );
  INV_X1 U34453 ( .A(n29982), .ZN(p_wishbone_bd_ram_n22913) );
  INV_X1 U34454 ( .A(n61237), .ZN(n29984) );
  INV_X1 U34455 ( .A(n29984), .ZN(p_wishbone_bd_ram_n22912) );
  INV_X1 U34456 ( .A(n61236), .ZN(n29986) );
  INV_X1 U34457 ( .A(n29986), .ZN(p_wishbone_bd_ram_n22911) );
  INV_X1 U34458 ( .A(n61235), .ZN(n29988) );
  INV_X1 U34459 ( .A(n29988), .ZN(p_wishbone_bd_ram_n22910) );
  INV_X1 U34460 ( .A(n61234), .ZN(n29990) );
  INV_X1 U34461 ( .A(n29990), .ZN(p_wishbone_bd_ram_n22909) );
  INV_X1 U34462 ( .A(n61233), .ZN(n29992) );
  INV_X1 U34463 ( .A(n29992), .ZN(p_wishbone_bd_ram_n22908) );
  INV_X1 U34464 ( .A(n61232), .ZN(n29994) );
  INV_X1 U34465 ( .A(n29994), .ZN(p_wishbone_bd_ram_n22907) );
  INV_X1 U34466 ( .A(n61231), .ZN(n29996) );
  INV_X1 U34467 ( .A(n29996), .ZN(p_wishbone_bd_ram_n22906) );
  INV_X1 U34468 ( .A(n61230), .ZN(n29998) );
  INV_X1 U34469 ( .A(n29998), .ZN(p_wishbone_bd_ram_n22905) );
  INV_X1 U34470 ( .A(n61229), .ZN(n30000) );
  INV_X1 U34471 ( .A(n30000), .ZN(p_wishbone_bd_ram_n22904) );
  INV_X1 U34472 ( .A(n61228), .ZN(n30002) );
  INV_X1 U34473 ( .A(n30002), .ZN(p_wishbone_bd_ram_n22903) );
  INV_X1 U34474 ( .A(n61227), .ZN(n30004) );
  INV_X1 U34475 ( .A(n30004), .ZN(p_wishbone_bd_ram_n22902) );
  INV_X1 U34476 ( .A(n61226), .ZN(n30006) );
  INV_X1 U34477 ( .A(n30006), .ZN(p_wishbone_bd_ram_n22901) );
  INV_X1 U34478 ( .A(n61225), .ZN(n30008) );
  INV_X1 U34479 ( .A(n30008), .ZN(p_wishbone_bd_ram_n22900) );
  INV_X1 U34480 ( .A(n61224), .ZN(n30010) );
  INV_X1 U34481 ( .A(n30010), .ZN(p_wishbone_bd_ram_n22899) );
  INV_X1 U34482 ( .A(n61223), .ZN(n30012) );
  INV_X1 U34483 ( .A(n30012), .ZN(p_wishbone_bd_ram_n22898) );
  INV_X1 U34484 ( .A(n61222), .ZN(n30014) );
  INV_X1 U34485 ( .A(n30014), .ZN(p_wishbone_bd_ram_n22897) );
  INV_X1 U34486 ( .A(n61221), .ZN(n30016) );
  INV_X1 U34487 ( .A(n30016), .ZN(p_wishbone_bd_ram_n22896) );
  INV_X1 U34488 ( .A(n61220), .ZN(n30018) );
  INV_X1 U34489 ( .A(n30018), .ZN(p_wishbone_bd_ram_n22895) );
  INV_X1 U34490 ( .A(n61219), .ZN(n30020) );
  INV_X1 U34491 ( .A(n30020), .ZN(p_wishbone_bd_ram_n22894) );
  INV_X1 U34492 ( .A(n61218), .ZN(n30022) );
  INV_X1 U34493 ( .A(n30022), .ZN(p_wishbone_bd_ram_n22893) );
  INV_X1 U34494 ( .A(n61217), .ZN(n30024) );
  INV_X1 U34495 ( .A(n30024), .ZN(p_wishbone_bd_ram_n22892) );
  INV_X1 U34496 ( .A(n61216), .ZN(n30026) );
  INV_X1 U34497 ( .A(n30026), .ZN(p_wishbone_bd_ram_n22891) );
  INV_X1 U34498 ( .A(n61215), .ZN(n30028) );
  INV_X1 U34499 ( .A(n30028), .ZN(p_wishbone_bd_ram_n22890) );
  INV_X1 U34500 ( .A(n61214), .ZN(n30030) );
  INV_X1 U34501 ( .A(n30030), .ZN(p_wishbone_bd_ram_n22889) );
  INV_X1 U34502 ( .A(n61213), .ZN(n30032) );
  INV_X1 U34503 ( .A(n30032), .ZN(p_wishbone_bd_ram_n22887) );
  INV_X1 U34504 ( .A(n61212), .ZN(n30034) );
  INV_X1 U34505 ( .A(n30034), .ZN(p_wishbone_bd_ram_n22885) );
  INV_X1 U34506 ( .A(n61211), .ZN(n30036) );
  INV_X1 U34507 ( .A(n30036), .ZN(p_wishbone_bd_ram_n22884) );
  INV_X1 U34508 ( .A(n61210), .ZN(n30038) );
  INV_X1 U34509 ( .A(n30038), .ZN(p_wishbone_bd_ram_n22882) );
  INV_X1 U34510 ( .A(n61209), .ZN(n30040) );
  INV_X1 U34511 ( .A(n30040), .ZN(p_wishbone_bd_ram_n22879) );
  INV_X1 U34512 ( .A(n61208), .ZN(n30042) );
  INV_X1 U34513 ( .A(n30042), .ZN(p_wishbone_bd_ram_n22877) );
  INV_X1 U34514 ( .A(n61207), .ZN(n30044) );
  INV_X1 U34515 ( .A(n30044), .ZN(p_wishbone_bd_ram_n22876) );
  INV_X1 U34516 ( .A(n61206), .ZN(n30046) );
  INV_X1 U34517 ( .A(n30046), .ZN(p_wishbone_bd_ram_n22874) );
  INV_X1 U34518 ( .A(n61205), .ZN(n30048) );
  INV_X1 U34519 ( .A(n30048), .ZN(p_wishbone_bd_ram_n22872) );
  INV_X1 U34520 ( .A(n61204), .ZN(n30050) );
  INV_X1 U34521 ( .A(n30050), .ZN(p_wishbone_bd_ram_n22871) );
  INV_X1 U34522 ( .A(n61203), .ZN(n30052) );
  INV_X1 U34523 ( .A(n30052), .ZN(p_wishbone_bd_ram_n22870) );
  INV_X1 U34524 ( .A(n61202), .ZN(n30054) );
  INV_X1 U34525 ( .A(n30054), .ZN(p_wishbone_bd_ram_n22869) );
  INV_X1 U34526 ( .A(n61201), .ZN(n30056) );
  INV_X1 U34527 ( .A(n30056), .ZN(p_wishbone_bd_ram_n22868) );
  INV_X1 U34528 ( .A(n61200), .ZN(n30058) );
  INV_X1 U34529 ( .A(n30058), .ZN(p_wishbone_bd_ram_n22867) );
  INV_X1 U34530 ( .A(n61199), .ZN(n30060) );
  INV_X1 U34531 ( .A(n30060), .ZN(p_wishbone_bd_ram_n22866) );
  INV_X1 U34532 ( .A(n61198), .ZN(n30062) );
  INV_X1 U34533 ( .A(n30062), .ZN(p_wishbone_bd_ram_n22865) );
  INV_X1 U34534 ( .A(n61197), .ZN(n30064) );
  INV_X1 U34535 ( .A(n30064), .ZN(p_wishbone_bd_ram_n22863) );
  INV_X1 U34536 ( .A(n61196), .ZN(n30066) );
  INV_X1 U34537 ( .A(n30066), .ZN(p_wishbone_bd_ram_n22861) );
  INV_X1 U34538 ( .A(n61195), .ZN(n30068) );
  INV_X1 U34539 ( .A(n30068), .ZN(p_wishbone_bd_ram_n22860) );
  INV_X1 U34540 ( .A(n61194), .ZN(n30070) );
  INV_X1 U34541 ( .A(n30070), .ZN(p_wishbone_bd_ram_n22858) );
  INV_X1 U34542 ( .A(n61193), .ZN(n30072) );
  INV_X1 U34543 ( .A(n30072), .ZN(p_wishbone_bd_ram_n22856) );
  INV_X1 U34544 ( .A(n61192), .ZN(n30074) );
  INV_X1 U34545 ( .A(n30074), .ZN(p_wishbone_bd_ram_n22855) );
  INV_X1 U34546 ( .A(n61191), .ZN(n30076) );
  INV_X1 U34547 ( .A(n30076), .ZN(p_wishbone_bd_ram_n22854) );
  INV_X1 U34548 ( .A(n61190), .ZN(n30078) );
  INV_X1 U34549 ( .A(n30078), .ZN(p_wishbone_bd_ram_n22853) );
  INV_X1 U34550 ( .A(n61189), .ZN(n30080) );
  INV_X1 U34551 ( .A(n30080), .ZN(p_wishbone_bd_ram_n22852) );
  INV_X1 U34552 ( .A(n61188), .ZN(n30082) );
  INV_X1 U34553 ( .A(n30082), .ZN(p_wishbone_bd_ram_n22851) );
  INV_X1 U34554 ( .A(n61187), .ZN(n30084) );
  INV_X1 U34555 ( .A(n30084), .ZN(p_wishbone_bd_ram_n22850) );
  INV_X1 U34556 ( .A(n61186), .ZN(n30086) );
  INV_X1 U34557 ( .A(n30086), .ZN(p_wishbone_bd_ram_n22849) );
  INV_X1 U34558 ( .A(n61185), .ZN(n30088) );
  INV_X1 U34559 ( .A(n30088), .ZN(p_wishbone_bd_ram_n22848) );
  INV_X1 U34560 ( .A(n61184), .ZN(n30090) );
  INV_X1 U34561 ( .A(n30090), .ZN(p_wishbone_bd_ram_n22847) );
  INV_X1 U34562 ( .A(n61183), .ZN(n30092) );
  INV_X1 U34563 ( .A(n30092), .ZN(p_wishbone_bd_ram_n22846) );
  INV_X1 U34564 ( .A(n61182), .ZN(n30094) );
  INV_X1 U34565 ( .A(n30094), .ZN(p_wishbone_bd_ram_n22845) );
  INV_X1 U34566 ( .A(n61181), .ZN(n30096) );
  INV_X1 U34567 ( .A(n30096), .ZN(p_wishbone_bd_ram_n22844) );
  INV_X1 U34568 ( .A(n61180), .ZN(n30098) );
  INV_X1 U34569 ( .A(n30098), .ZN(p_wishbone_bd_ram_n22843) );
  INV_X1 U34570 ( .A(n61179), .ZN(n30100) );
  INV_X1 U34571 ( .A(n30100), .ZN(p_wishbone_bd_ram_n22842) );
  INV_X1 U34572 ( .A(n61178), .ZN(n30102) );
  INV_X1 U34573 ( .A(n30102), .ZN(p_wishbone_bd_ram_n22841) );
  INV_X1 U34574 ( .A(n61177), .ZN(n30104) );
  INV_X1 U34575 ( .A(n30104), .ZN(p_wishbone_bd_ram_n22840) );
  INV_X1 U34576 ( .A(n61176), .ZN(n30106) );
  INV_X1 U34577 ( .A(n30106), .ZN(p_wishbone_bd_ram_n22839) );
  INV_X1 U34578 ( .A(n61175), .ZN(n30108) );
  INV_X1 U34579 ( .A(n30108), .ZN(p_wishbone_bd_ram_n22838) );
  INV_X1 U34580 ( .A(n61174), .ZN(n30110) );
  INV_X1 U34581 ( .A(n30110), .ZN(p_wishbone_bd_ram_n22837) );
  INV_X1 U34582 ( .A(n61173), .ZN(n30112) );
  INV_X1 U34583 ( .A(n30112), .ZN(p_wishbone_bd_ram_n22836) );
  INV_X1 U34584 ( .A(n61172), .ZN(n30114) );
  INV_X1 U34585 ( .A(n30114), .ZN(p_wishbone_bd_ram_n22835) );
  INV_X1 U34586 ( .A(n61171), .ZN(n30116) );
  INV_X1 U34587 ( .A(n30116), .ZN(p_wishbone_bd_ram_n22834) );
  INV_X1 U34588 ( .A(n61170), .ZN(n30118) );
  INV_X1 U34589 ( .A(n30118), .ZN(p_wishbone_bd_ram_n22833) );
  INV_X1 U34590 ( .A(n61169), .ZN(n30120) );
  INV_X1 U34591 ( .A(n30120), .ZN(p_wishbone_bd_ram_n22832) );
  INV_X1 U34592 ( .A(n61168), .ZN(n30122) );
  INV_X1 U34593 ( .A(n30122), .ZN(p_wishbone_bd_ram_n22831) );
  INV_X1 U34594 ( .A(n61167), .ZN(n30124) );
  INV_X1 U34595 ( .A(n30124), .ZN(p_wishbone_bd_ram_n22830) );
  INV_X1 U34596 ( .A(n61166), .ZN(n30126) );
  INV_X1 U34597 ( .A(n30126), .ZN(p_wishbone_bd_ram_n22829) );
  INV_X1 U34598 ( .A(n61165), .ZN(n30128) );
  INV_X1 U34599 ( .A(n30128), .ZN(p_wishbone_bd_ram_n22828) );
  INV_X1 U34600 ( .A(n61164), .ZN(n30130) );
  INV_X1 U34601 ( .A(n30130), .ZN(p_wishbone_bd_ram_n22827) );
  INV_X1 U34602 ( .A(n61163), .ZN(n30132) );
  INV_X1 U34603 ( .A(n30132), .ZN(p_wishbone_bd_ram_n22826) );
  INV_X1 U34604 ( .A(n61162), .ZN(n30134) );
  INV_X1 U34605 ( .A(n30134), .ZN(p_wishbone_bd_ram_n22825) );
  INV_X1 U34606 ( .A(n61161), .ZN(n30136) );
  INV_X1 U34607 ( .A(n30136), .ZN(p_wishbone_bd_ram_n22823) );
  INV_X1 U34608 ( .A(n61160), .ZN(n30138) );
  INV_X1 U34609 ( .A(n30138), .ZN(p_wishbone_bd_ram_n22821) );
  INV_X1 U34610 ( .A(n61159), .ZN(n30140) );
  INV_X1 U34611 ( .A(n30140), .ZN(p_wishbone_bd_ram_n22820) );
  INV_X1 U34612 ( .A(n61158), .ZN(n30142) );
  INV_X1 U34613 ( .A(n30142), .ZN(p_wishbone_bd_ram_n22818) );
  INV_X1 U34614 ( .A(n61157), .ZN(n30144) );
  INV_X1 U34615 ( .A(n30144), .ZN(p_wishbone_bd_ram_n22816) );
  INV_X1 U34616 ( .A(n61156), .ZN(n30146) );
  INV_X1 U34617 ( .A(n30146), .ZN(p_wishbone_bd_ram_n22815) );
  INV_X1 U34618 ( .A(n61155), .ZN(n30148) );
  INV_X1 U34619 ( .A(n30148), .ZN(p_wishbone_bd_ram_n22814) );
  INV_X1 U34620 ( .A(n61154), .ZN(n30150) );
  INV_X1 U34621 ( .A(n30150), .ZN(p_wishbone_bd_ram_n22813) );
  INV_X1 U34622 ( .A(n61153), .ZN(n30152) );
  INV_X1 U34623 ( .A(n30152), .ZN(p_wishbone_bd_ram_n22812) );
  INV_X1 U34624 ( .A(n61152), .ZN(n30154) );
  INV_X1 U34625 ( .A(n30154), .ZN(p_wishbone_bd_ram_n22811) );
  INV_X1 U34626 ( .A(n61151), .ZN(n30156) );
  INV_X1 U34627 ( .A(n30156), .ZN(p_wishbone_bd_ram_n22810) );
  INV_X1 U34628 ( .A(n61150), .ZN(n30158) );
  INV_X1 U34629 ( .A(n30158), .ZN(p_wishbone_bd_ram_n22809) );
  INV_X1 U34630 ( .A(n61149), .ZN(n30160) );
  INV_X1 U34631 ( .A(n30160), .ZN(p_wishbone_bd_ram_n22808) );
  INV_X1 U34632 ( .A(n61148), .ZN(n30162) );
  INV_X1 U34633 ( .A(n30162), .ZN(p_wishbone_bd_ram_n22807) );
  INV_X1 U34634 ( .A(n61147), .ZN(n30164) );
  INV_X1 U34635 ( .A(n30164), .ZN(p_wishbone_bd_ram_n22806) );
  INV_X1 U34636 ( .A(n61146), .ZN(n30166) );
  INV_X1 U34637 ( .A(n30166), .ZN(p_wishbone_bd_ram_n22805) );
  INV_X1 U34638 ( .A(n61145), .ZN(n30168) );
  INV_X1 U34639 ( .A(n30168), .ZN(p_wishbone_bd_ram_n22804) );
  INV_X1 U34640 ( .A(n61144), .ZN(n30170) );
  INV_X1 U34641 ( .A(n30170), .ZN(p_wishbone_bd_ram_n22803) );
  INV_X1 U34642 ( .A(n61143), .ZN(n30172) );
  INV_X1 U34643 ( .A(n30172), .ZN(p_wishbone_bd_ram_n22802) );
  INV_X1 U34644 ( .A(n61142), .ZN(n30174) );
  INV_X1 U34645 ( .A(n30174), .ZN(p_wishbone_bd_ram_n22801) );
  INV_X1 U34646 ( .A(n61141), .ZN(n30176) );
  INV_X1 U34647 ( .A(n30176), .ZN(p_wishbone_bd_ram_n22800) );
  INV_X1 U34648 ( .A(n61140), .ZN(n30178) );
  INV_X1 U34649 ( .A(n30178), .ZN(p_wishbone_bd_ram_n22799) );
  INV_X1 U34650 ( .A(n61139), .ZN(n30180) );
  INV_X1 U34651 ( .A(n30180), .ZN(p_wishbone_bd_ram_n22798) );
  INV_X1 U34652 ( .A(n61138), .ZN(n30182) );
  INV_X1 U34653 ( .A(n30182), .ZN(p_wishbone_bd_ram_n22797) );
  INV_X1 U34654 ( .A(n61137), .ZN(n30184) );
  INV_X1 U34655 ( .A(n30184), .ZN(p_wishbone_bd_ram_n22796) );
  INV_X1 U34656 ( .A(n61136), .ZN(n30186) );
  INV_X1 U34657 ( .A(n30186), .ZN(p_wishbone_bd_ram_n22795) );
  INV_X1 U34658 ( .A(n61135), .ZN(n30188) );
  INV_X1 U34659 ( .A(n30188), .ZN(p_wishbone_bd_ram_n22794) );
  INV_X1 U34660 ( .A(n61134), .ZN(n30190) );
  INV_X1 U34661 ( .A(n30190), .ZN(p_wishbone_bd_ram_n22793) );
  INV_X1 U34662 ( .A(n61133), .ZN(n30192) );
  INV_X1 U34663 ( .A(n30192), .ZN(p_wishbone_bd_ram_n22792) );
  INV_X1 U34664 ( .A(n61132), .ZN(n30194) );
  INV_X1 U34665 ( .A(n30194), .ZN(p_wishbone_bd_ram_n22791) );
  INV_X1 U34666 ( .A(n61131), .ZN(n30196) );
  INV_X1 U34667 ( .A(n30196), .ZN(p_wishbone_bd_ram_n22790) );
  INV_X1 U34668 ( .A(n61130), .ZN(n30198) );
  INV_X1 U34669 ( .A(n30198), .ZN(p_wishbone_bd_ram_n22789) );
  INV_X1 U34670 ( .A(n61129), .ZN(n30200) );
  INV_X1 U34671 ( .A(n30200), .ZN(p_wishbone_bd_ram_n22788) );
  INV_X1 U34672 ( .A(n61128), .ZN(n30202) );
  INV_X1 U34673 ( .A(n30202), .ZN(p_wishbone_bd_ram_n22787) );
  INV_X1 U34674 ( .A(n61127), .ZN(n30204) );
  INV_X1 U34675 ( .A(n30204), .ZN(p_wishbone_bd_ram_n22786) );
  INV_X1 U34676 ( .A(n61126), .ZN(n30206) );
  INV_X1 U34677 ( .A(n30206), .ZN(p_wishbone_bd_ram_n22785) );
  INV_X1 U34678 ( .A(n61125), .ZN(n30208) );
  INV_X1 U34679 ( .A(n30208), .ZN(p_wishbone_bd_ram_n22784) );
  INV_X1 U34680 ( .A(n61124), .ZN(n30210) );
  INV_X1 U34681 ( .A(n30210), .ZN(p_wishbone_bd_ram_n22783) );
  INV_X1 U34682 ( .A(n61123), .ZN(n30212) );
  INV_X1 U34683 ( .A(n30212), .ZN(p_wishbone_bd_ram_n22782) );
  INV_X1 U34684 ( .A(n61122), .ZN(n30214) );
  INV_X1 U34685 ( .A(n30214), .ZN(p_wishbone_bd_ram_n22781) );
  INV_X1 U34686 ( .A(n61121), .ZN(n30216) );
  INV_X1 U34687 ( .A(n30216), .ZN(p_wishbone_bd_ram_n22780) );
  INV_X1 U34688 ( .A(n61120), .ZN(n30218) );
  INV_X1 U34689 ( .A(n30218), .ZN(p_wishbone_bd_ram_n22779) );
  INV_X1 U34690 ( .A(n61119), .ZN(n30220) );
  INV_X1 U34691 ( .A(n30220), .ZN(p_wishbone_bd_ram_n22778) );
  INV_X1 U34692 ( .A(n61118), .ZN(n30222) );
  INV_X1 U34693 ( .A(n30222), .ZN(p_wishbone_bd_ram_n22777) );
  INV_X1 U34694 ( .A(n61117), .ZN(n30224) );
  INV_X1 U34695 ( .A(n30224), .ZN(p_wishbone_bd_ram_n22776) );
  INV_X1 U34696 ( .A(n61116), .ZN(n30226) );
  INV_X1 U34697 ( .A(n30226), .ZN(p_wishbone_bd_ram_n22775) );
  INV_X1 U34698 ( .A(n61115), .ZN(n30228) );
  INV_X1 U34699 ( .A(n30228), .ZN(p_wishbone_bd_ram_n22774) );
  INV_X1 U34700 ( .A(n61114), .ZN(n30230) );
  INV_X1 U34701 ( .A(n30230), .ZN(p_wishbone_bd_ram_n22773) );
  INV_X1 U34702 ( .A(n61113), .ZN(n30232) );
  INV_X1 U34703 ( .A(n30232), .ZN(p_wishbone_bd_ram_n22772) );
  INV_X1 U34704 ( .A(n61112), .ZN(n30234) );
  INV_X1 U34705 ( .A(n30234), .ZN(p_wishbone_bd_ram_n22771) );
  INV_X1 U34706 ( .A(n61111), .ZN(n30236) );
  INV_X1 U34707 ( .A(n30236), .ZN(p_wishbone_bd_ram_n22770) );
  INV_X1 U34708 ( .A(n61110), .ZN(n30238) );
  INV_X1 U34709 ( .A(n30238), .ZN(p_wishbone_bd_ram_n22769) );
  INV_X1 U34710 ( .A(n61109), .ZN(n30240) );
  INV_X1 U34711 ( .A(n30240), .ZN(p_wishbone_bd_ram_n22768) );
  INV_X1 U34712 ( .A(n61108), .ZN(n30242) );
  INV_X1 U34713 ( .A(n30242), .ZN(p_wishbone_bd_ram_n22767) );
  INV_X1 U34714 ( .A(n61107), .ZN(n30244) );
  INV_X1 U34715 ( .A(n30244), .ZN(p_wishbone_bd_ram_n22766) );
  INV_X1 U34716 ( .A(n61106), .ZN(n30246) );
  INV_X1 U34717 ( .A(n30246), .ZN(p_wishbone_bd_ram_n22765) );
  INV_X1 U34718 ( .A(n61105), .ZN(n30248) );
  INV_X1 U34719 ( .A(n30248), .ZN(p_wishbone_bd_ram_n22764) );
  INV_X1 U34720 ( .A(n61104), .ZN(n30250) );
  INV_X1 U34721 ( .A(n30250), .ZN(p_wishbone_bd_ram_n22763) );
  INV_X1 U34722 ( .A(n61103), .ZN(n30252) );
  INV_X1 U34723 ( .A(n30252), .ZN(p_wishbone_bd_ram_n22762) );
  INV_X1 U34724 ( .A(n61102), .ZN(n30254) );
  INV_X1 U34725 ( .A(n30254), .ZN(p_wishbone_bd_ram_n22761) );
  INV_X1 U34726 ( .A(n61101), .ZN(n30256) );
  INV_X1 U34727 ( .A(n30256), .ZN(p_wishbone_bd_ram_n22759) );
  INV_X1 U34728 ( .A(n61100), .ZN(n30258) );
  INV_X1 U34729 ( .A(n30258), .ZN(p_wishbone_bd_ram_n22757) );
  INV_X1 U34730 ( .A(n61099), .ZN(n30260) );
  INV_X1 U34731 ( .A(n30260), .ZN(p_wishbone_bd_ram_n22756) );
  INV_X1 U34732 ( .A(n61098), .ZN(n30262) );
  INV_X1 U34733 ( .A(n30262), .ZN(p_wishbone_bd_ram_n22754) );
  INV_X1 U34734 ( .A(n61097), .ZN(n30264) );
  INV_X1 U34735 ( .A(n30264), .ZN(p_wishbone_bd_ram_n22752) );
  INV_X1 U34736 ( .A(n61096), .ZN(n30266) );
  INV_X1 U34737 ( .A(n30266), .ZN(p_wishbone_bd_ram_n22751) );
  INV_X1 U34738 ( .A(n61095), .ZN(n30268) );
  INV_X1 U34739 ( .A(n30268), .ZN(p_wishbone_bd_ram_n22750) );
  INV_X1 U34740 ( .A(n61094), .ZN(n30270) );
  INV_X1 U34741 ( .A(n30270), .ZN(p_wishbone_bd_ram_n22749) );
  INV_X1 U34742 ( .A(n61093), .ZN(n30272) );
  INV_X1 U34743 ( .A(n30272), .ZN(p_wishbone_bd_ram_n22748) );
  INV_X1 U34744 ( .A(n61092), .ZN(n30274) );
  INV_X1 U34745 ( .A(n30274), .ZN(p_wishbone_bd_ram_n22747) );
  INV_X1 U34746 ( .A(n61091), .ZN(n30276) );
  INV_X1 U34747 ( .A(n30276), .ZN(p_wishbone_bd_ram_n22746) );
  INV_X1 U34748 ( .A(n61090), .ZN(n30278) );
  INV_X1 U34749 ( .A(n30278), .ZN(p_wishbone_bd_ram_n22745) );
  INV_X1 U34750 ( .A(n61089), .ZN(n30280) );
  INV_X1 U34751 ( .A(n30280), .ZN(p_wishbone_bd_ram_n22744) );
  INV_X1 U34752 ( .A(n61088), .ZN(n30282) );
  INV_X1 U34753 ( .A(n30282), .ZN(p_wishbone_bd_ram_n22743) );
  INV_X1 U34754 ( .A(n61087), .ZN(n30284) );
  INV_X1 U34755 ( .A(n30284), .ZN(p_wishbone_bd_ram_n22742) );
  INV_X1 U34756 ( .A(n61086), .ZN(n30286) );
  INV_X1 U34757 ( .A(n30286), .ZN(p_wishbone_bd_ram_n22741) );
  INV_X1 U34758 ( .A(n61085), .ZN(n30288) );
  INV_X1 U34759 ( .A(n30288), .ZN(p_wishbone_bd_ram_n22740) );
  INV_X1 U34760 ( .A(n61084), .ZN(n30290) );
  INV_X1 U34761 ( .A(n30290), .ZN(p_wishbone_bd_ram_n22739) );
  INV_X1 U34762 ( .A(n61083), .ZN(n30292) );
  INV_X1 U34763 ( .A(n30292), .ZN(p_wishbone_bd_ram_n22738) );
  INV_X1 U34764 ( .A(n61082), .ZN(n30294) );
  INV_X1 U34765 ( .A(n30294), .ZN(p_wishbone_bd_ram_n22737) );
  INV_X1 U34766 ( .A(n61081), .ZN(n30296) );
  INV_X1 U34767 ( .A(n30296), .ZN(p_wishbone_bd_ram_n22735) );
  INV_X1 U34768 ( .A(n61080), .ZN(n30298) );
  INV_X1 U34769 ( .A(n30298), .ZN(p_wishbone_bd_ram_n22733) );
  INV_X1 U34770 ( .A(n61079), .ZN(n30300) );
  INV_X1 U34771 ( .A(n30300), .ZN(p_wishbone_bd_ram_n22732) );
  INV_X1 U34772 ( .A(n61078), .ZN(n30302) );
  INV_X1 U34773 ( .A(n30302), .ZN(p_wishbone_bd_ram_n22730) );
  INV_X1 U34774 ( .A(n61077), .ZN(n30304) );
  INV_X1 U34775 ( .A(n30304), .ZN(p_wishbone_bd_ram_n22728) );
  INV_X1 U34776 ( .A(n61076), .ZN(n30306) );
  INV_X1 U34777 ( .A(n30306), .ZN(p_wishbone_bd_ram_n22727) );
  INV_X1 U34778 ( .A(n61075), .ZN(n30308) );
  INV_X1 U34779 ( .A(n30308), .ZN(p_wishbone_bd_ram_n22726) );
  INV_X1 U34780 ( .A(n61074), .ZN(n30310) );
  INV_X1 U34781 ( .A(n30310), .ZN(p_wishbone_bd_ram_n22725) );
  INV_X1 U34782 ( .A(n61073), .ZN(n30312) );
  INV_X1 U34783 ( .A(n30312), .ZN(p_wishbone_bd_ram_n22724) );
  INV_X1 U34784 ( .A(n61072), .ZN(n30314) );
  INV_X1 U34785 ( .A(n30314), .ZN(p_wishbone_bd_ram_n22723) );
  INV_X1 U34786 ( .A(n61071), .ZN(n30316) );
  INV_X1 U34787 ( .A(n30316), .ZN(p_wishbone_bd_ram_n22722) );
  INV_X1 U34788 ( .A(n61070), .ZN(n30318) );
  INV_X1 U34789 ( .A(n30318), .ZN(p_wishbone_bd_ram_n22721) );
  INV_X1 U34790 ( .A(n61069), .ZN(n30320) );
  INV_X1 U34791 ( .A(n30320), .ZN(p_wishbone_bd_ram_n22720) );
  INV_X1 U34792 ( .A(n61068), .ZN(n30322) );
  INV_X1 U34793 ( .A(n30322), .ZN(p_wishbone_bd_ram_n22719) );
  INV_X1 U34794 ( .A(n61067), .ZN(n30324) );
  INV_X1 U34795 ( .A(n30324), .ZN(p_wishbone_bd_ram_n22718) );
  INV_X1 U34796 ( .A(n61066), .ZN(n30326) );
  INV_X1 U34797 ( .A(n30326), .ZN(p_wishbone_bd_ram_n22717) );
  INV_X1 U34798 ( .A(n61065), .ZN(n30328) );
  INV_X1 U34799 ( .A(n30328), .ZN(p_wishbone_bd_ram_n22716) );
  INV_X1 U34800 ( .A(n61064), .ZN(n30330) );
  INV_X1 U34801 ( .A(n30330), .ZN(p_wishbone_bd_ram_n22715) );
  INV_X1 U34802 ( .A(n61063), .ZN(n30332) );
  INV_X1 U34803 ( .A(n30332), .ZN(p_wishbone_bd_ram_n22714) );
  INV_X1 U34804 ( .A(n61062), .ZN(n30334) );
  INV_X1 U34805 ( .A(n30334), .ZN(p_wishbone_bd_ram_n22713) );
  INV_X1 U34806 ( .A(n61061), .ZN(n30336) );
  INV_X1 U34807 ( .A(n30336), .ZN(p_wishbone_bd_ram_n22712) );
  INV_X1 U34808 ( .A(n61060), .ZN(n30338) );
  INV_X1 U34809 ( .A(n30338), .ZN(p_wishbone_bd_ram_n22711) );
  INV_X1 U34810 ( .A(n61059), .ZN(n30340) );
  INV_X1 U34811 ( .A(n30340), .ZN(p_wishbone_bd_ram_n22710) );
  INV_X1 U34812 ( .A(n61058), .ZN(n30342) );
  INV_X1 U34813 ( .A(n30342), .ZN(p_wishbone_bd_ram_n22709) );
  INV_X1 U34814 ( .A(n61057), .ZN(n30344) );
  INV_X1 U34815 ( .A(n30344), .ZN(p_wishbone_bd_ram_n22708) );
  INV_X1 U34816 ( .A(n61056), .ZN(n30346) );
  INV_X1 U34817 ( .A(n30346), .ZN(p_wishbone_bd_ram_n22707) );
  INV_X1 U34818 ( .A(n61055), .ZN(n30348) );
  INV_X1 U34819 ( .A(n30348), .ZN(p_wishbone_bd_ram_n22706) );
  INV_X1 U34820 ( .A(n61054), .ZN(n30350) );
  INV_X1 U34821 ( .A(n30350), .ZN(p_wishbone_bd_ram_n22705) );
  INV_X1 U34822 ( .A(n61053), .ZN(n30352) );
  INV_X1 U34823 ( .A(n30352), .ZN(p_wishbone_bd_ram_n22704) );
  INV_X1 U34824 ( .A(n61052), .ZN(n30354) );
  INV_X1 U34825 ( .A(n30354), .ZN(p_wishbone_bd_ram_n22703) );
  INV_X1 U34826 ( .A(n61051), .ZN(n30356) );
  INV_X1 U34827 ( .A(n30356), .ZN(p_wishbone_bd_ram_n22702) );
  INV_X1 U34828 ( .A(n61050), .ZN(n30358) );
  INV_X1 U34829 ( .A(n30358), .ZN(p_wishbone_bd_ram_n22701) );
  INV_X1 U34830 ( .A(n61049), .ZN(n30360) );
  INV_X1 U34831 ( .A(n30360), .ZN(p_wishbone_bd_ram_n22700) );
  INV_X1 U34832 ( .A(n61048), .ZN(n30362) );
  INV_X1 U34833 ( .A(n30362), .ZN(p_wishbone_bd_ram_n22699) );
  INV_X1 U34834 ( .A(n61047), .ZN(n30364) );
  INV_X1 U34835 ( .A(n30364), .ZN(p_wishbone_bd_ram_n22698) );
  INV_X1 U34836 ( .A(n61046), .ZN(n30366) );
  INV_X1 U34837 ( .A(n30366), .ZN(p_wishbone_bd_ram_n22697) );
  INV_X1 U34838 ( .A(n61045), .ZN(n30368) );
  INV_X1 U34839 ( .A(n30368), .ZN(p_wishbone_bd_ram_n22696) );
  INV_X1 U34840 ( .A(n61044), .ZN(n30370) );
  INV_X1 U34841 ( .A(n30370), .ZN(p_wishbone_bd_ram_n22695) );
  INV_X1 U34842 ( .A(n61043), .ZN(n30372) );
  INV_X1 U34843 ( .A(n30372), .ZN(p_wishbone_bd_ram_n22694) );
  INV_X1 U34844 ( .A(n61042), .ZN(n30374) );
  INV_X1 U34845 ( .A(n30374), .ZN(p_wishbone_bd_ram_n22693) );
  INV_X1 U34846 ( .A(n61041), .ZN(n30376) );
  INV_X1 U34847 ( .A(n30376), .ZN(p_wishbone_bd_ram_n22692) );
  INV_X1 U34848 ( .A(n61040), .ZN(n30378) );
  INV_X1 U34849 ( .A(n30378), .ZN(p_wishbone_bd_ram_n22691) );
  INV_X1 U34850 ( .A(n61039), .ZN(n30380) );
  INV_X1 U34851 ( .A(n30380), .ZN(p_wishbone_bd_ram_n22690) );
  INV_X1 U34852 ( .A(n61038), .ZN(n30382) );
  INV_X1 U34853 ( .A(n30382), .ZN(p_wishbone_bd_ram_n22689) );
  INV_X1 U34854 ( .A(n61037), .ZN(n30384) );
  INV_X1 U34855 ( .A(n30384), .ZN(p_wishbone_bd_ram_n22688) );
  INV_X1 U34856 ( .A(n61036), .ZN(n30386) );
  INV_X1 U34857 ( .A(n30386), .ZN(p_wishbone_bd_ram_n22687) );
  INV_X1 U34858 ( .A(n61035), .ZN(n30388) );
  INV_X1 U34859 ( .A(n30388), .ZN(p_wishbone_bd_ram_n22686) );
  INV_X1 U34860 ( .A(n61034), .ZN(n30390) );
  INV_X1 U34861 ( .A(n30390), .ZN(p_wishbone_bd_ram_n22685) );
  INV_X1 U34862 ( .A(n61033), .ZN(n30392) );
  INV_X1 U34863 ( .A(n30392), .ZN(p_wishbone_bd_ram_n22684) );
  INV_X1 U34864 ( .A(n61032), .ZN(n30394) );
  INV_X1 U34865 ( .A(n30394), .ZN(p_wishbone_bd_ram_n22683) );
  INV_X1 U34866 ( .A(n61031), .ZN(n30396) );
  INV_X1 U34867 ( .A(n30396), .ZN(p_wishbone_bd_ram_n22682) );
  INV_X1 U34868 ( .A(n61030), .ZN(n30398) );
  INV_X1 U34869 ( .A(n30398), .ZN(p_wishbone_bd_ram_n22681) );
  INV_X1 U34870 ( .A(n61029), .ZN(n30400) );
  INV_X1 U34871 ( .A(n30400), .ZN(p_wishbone_bd_ram_n22680) );
  INV_X1 U34872 ( .A(n61028), .ZN(n30402) );
  INV_X1 U34873 ( .A(n30402), .ZN(p_wishbone_bd_ram_n22679) );
  INV_X1 U34874 ( .A(n61027), .ZN(n30404) );
  INV_X1 U34875 ( .A(n30404), .ZN(p_wishbone_bd_ram_n22678) );
  INV_X1 U34876 ( .A(n61026), .ZN(n30406) );
  INV_X1 U34877 ( .A(n30406), .ZN(p_wishbone_bd_ram_n22677) );
  INV_X1 U34878 ( .A(n61025), .ZN(n30408) );
  INV_X1 U34879 ( .A(n30408), .ZN(p_wishbone_bd_ram_n22676) );
  INV_X1 U34880 ( .A(n61024), .ZN(n30410) );
  INV_X1 U34881 ( .A(n30410), .ZN(p_wishbone_bd_ram_n22675) );
  INV_X1 U34882 ( .A(n61023), .ZN(n30412) );
  INV_X1 U34883 ( .A(n30412), .ZN(p_wishbone_bd_ram_n22674) );
  INV_X1 U34884 ( .A(n61022), .ZN(n30414) );
  INV_X1 U34885 ( .A(n30414), .ZN(p_wishbone_bd_ram_n22673) );
  INV_X1 U34886 ( .A(n61021), .ZN(n30416) );
  INV_X1 U34887 ( .A(n30416), .ZN(p_wishbone_bd_ram_n22672) );
  INV_X1 U34888 ( .A(n61020), .ZN(n30418) );
  INV_X1 U34889 ( .A(n30418), .ZN(p_wishbone_bd_ram_n22671) );
  INV_X1 U34890 ( .A(n61019), .ZN(n30420) );
  INV_X1 U34891 ( .A(n30420), .ZN(p_wishbone_bd_ram_n22670) );
  INV_X1 U34892 ( .A(n61018), .ZN(n30422) );
  INV_X1 U34893 ( .A(n30422), .ZN(p_wishbone_bd_ram_n22669) );
  INV_X1 U34894 ( .A(n61017), .ZN(n30424) );
  INV_X1 U34895 ( .A(n30424), .ZN(p_wishbone_bd_ram_n22668) );
  INV_X1 U34896 ( .A(n61016), .ZN(n30426) );
  INV_X1 U34897 ( .A(n30426), .ZN(p_wishbone_bd_ram_n22667) );
  INV_X1 U34898 ( .A(n61015), .ZN(n30428) );
  INV_X1 U34899 ( .A(n30428), .ZN(p_wishbone_bd_ram_n22666) );
  INV_X1 U34900 ( .A(n61014), .ZN(n30430) );
  INV_X1 U34901 ( .A(n30430), .ZN(p_wishbone_bd_ram_n22665) );
  INV_X1 U34902 ( .A(n61013), .ZN(n30432) );
  INV_X1 U34903 ( .A(n30432), .ZN(p_wishbone_bd_ram_n22663) );
  INV_X1 U34904 ( .A(n61012), .ZN(n30434) );
  INV_X1 U34905 ( .A(n30434), .ZN(p_wishbone_bd_ram_n22661) );
  INV_X1 U34906 ( .A(n61011), .ZN(n30436) );
  INV_X1 U34907 ( .A(n30436), .ZN(p_wishbone_bd_ram_n22660) );
  INV_X1 U34908 ( .A(n61010), .ZN(n30438) );
  INV_X1 U34909 ( .A(n30438), .ZN(p_wishbone_bd_ram_n22658) );
  INV_X1 U34910 ( .A(n61009), .ZN(n30440) );
  INV_X1 U34911 ( .A(n30440), .ZN(p_wishbone_bd_ram_n22656) );
  INV_X1 U34912 ( .A(n61008), .ZN(n30442) );
  INV_X1 U34913 ( .A(n30442), .ZN(p_wishbone_bd_ram_n22655) );
  INV_X1 U34914 ( .A(n61007), .ZN(n30444) );
  INV_X1 U34915 ( .A(n30444), .ZN(p_wishbone_bd_ram_n22654) );
  INV_X1 U34916 ( .A(n61006), .ZN(n30446) );
  INV_X1 U34917 ( .A(n30446), .ZN(p_wishbone_bd_ram_n22653) );
  INV_X1 U34918 ( .A(n61005), .ZN(n30448) );
  INV_X1 U34919 ( .A(n30448), .ZN(p_wishbone_bd_ram_n22652) );
  INV_X1 U34920 ( .A(n61004), .ZN(n30450) );
  INV_X1 U34921 ( .A(n30450), .ZN(p_wishbone_bd_ram_n22651) );
  INV_X1 U34922 ( .A(n61003), .ZN(n30452) );
  INV_X1 U34923 ( .A(n30452), .ZN(p_wishbone_bd_ram_n22650) );
  INV_X1 U34924 ( .A(n61002), .ZN(n30454) );
  INV_X1 U34925 ( .A(n30454), .ZN(p_wishbone_bd_ram_n22649) );
  INV_X1 U34926 ( .A(n61001), .ZN(n30456) );
  INV_X1 U34927 ( .A(n30456), .ZN(p_wishbone_bd_ram_n22648) );
  INV_X1 U34928 ( .A(n61000), .ZN(n30458) );
  INV_X1 U34929 ( .A(n30458), .ZN(p_wishbone_bd_ram_n22647) );
  INV_X1 U34930 ( .A(n60999), .ZN(n30460) );
  INV_X1 U34931 ( .A(n30460), .ZN(p_wishbone_bd_ram_n22646) );
  INV_X1 U34932 ( .A(n60998), .ZN(n30462) );
  INV_X1 U34933 ( .A(n30462), .ZN(p_wishbone_bd_ram_n22645) );
  INV_X1 U34934 ( .A(n60997), .ZN(n30464) );
  INV_X1 U34935 ( .A(n30464), .ZN(p_wishbone_bd_ram_n22644) );
  INV_X1 U34936 ( .A(n60996), .ZN(n30466) );
  INV_X1 U34937 ( .A(n30466), .ZN(p_wishbone_bd_ram_n22643) );
  INV_X1 U34938 ( .A(n60995), .ZN(n30468) );
  INV_X1 U34939 ( .A(n30468), .ZN(p_wishbone_bd_ram_n22642) );
  INV_X1 U34940 ( .A(n60994), .ZN(n30470) );
  INV_X1 U34941 ( .A(n30470), .ZN(p_wishbone_bd_ram_n22641) );
  INV_X1 U34942 ( .A(n60993), .ZN(n30472) );
  INV_X1 U34943 ( .A(n30472), .ZN(p_wishbone_bd_ram_n22639) );
  INV_X1 U34944 ( .A(n60992), .ZN(n30474) );
  INV_X1 U34945 ( .A(n30474), .ZN(p_wishbone_bd_ram_n22637) );
  INV_X1 U34946 ( .A(n60991), .ZN(n30476) );
  INV_X1 U34947 ( .A(n30476), .ZN(p_wishbone_bd_ram_n22636) );
  INV_X1 U34948 ( .A(n60990), .ZN(n30478) );
  INV_X1 U34949 ( .A(n30478), .ZN(p_wishbone_bd_ram_n22634) );
  INV_X1 U34950 ( .A(n60989), .ZN(n30480) );
  INV_X1 U34951 ( .A(n30480), .ZN(p_wishbone_bd_ram_n22632) );
  INV_X1 U34952 ( .A(n60988), .ZN(n30482) );
  INV_X1 U34953 ( .A(n30482), .ZN(p_wishbone_bd_ram_n22631) );
  INV_X1 U34954 ( .A(n60987), .ZN(n30484) );
  INV_X1 U34955 ( .A(n30484), .ZN(p_wishbone_bd_ram_n22630) );
  INV_X1 U34956 ( .A(n60986), .ZN(n30486) );
  INV_X1 U34957 ( .A(n30486), .ZN(p_wishbone_bd_ram_n22629) );
  INV_X1 U34958 ( .A(n60985), .ZN(n30488) );
  INV_X1 U34959 ( .A(n30488), .ZN(p_wishbone_bd_ram_n22628) );
  INV_X1 U34960 ( .A(n60984), .ZN(n30490) );
  INV_X1 U34961 ( .A(n30490), .ZN(p_wishbone_bd_ram_n22627) );
  INV_X1 U34962 ( .A(n60983), .ZN(n30492) );
  INV_X1 U34963 ( .A(n30492), .ZN(p_wishbone_bd_ram_n22626) );
  INV_X1 U34964 ( .A(n60982), .ZN(n30494) );
  INV_X1 U34965 ( .A(n30494), .ZN(p_wishbone_bd_ram_n22625) );
  INV_X1 U34966 ( .A(n60981), .ZN(n30496) );
  INV_X1 U34967 ( .A(n30496), .ZN(p_wishbone_bd_ram_n22624) );
  INV_X1 U34968 ( .A(n60980), .ZN(n30498) );
  INV_X1 U34969 ( .A(n30498), .ZN(p_wishbone_bd_ram_n22623) );
  INV_X1 U34970 ( .A(n60979), .ZN(n30500) );
  INV_X1 U34971 ( .A(n30500), .ZN(p_wishbone_bd_ram_n22622) );
  INV_X1 U34972 ( .A(n60978), .ZN(n30502) );
  INV_X1 U34973 ( .A(n30502), .ZN(p_wishbone_bd_ram_n22621) );
  INV_X1 U34974 ( .A(n60977), .ZN(n30504) );
  INV_X1 U34975 ( .A(n30504), .ZN(p_wishbone_bd_ram_n22620) );
  INV_X1 U34976 ( .A(n60976), .ZN(n30506) );
  INV_X1 U34977 ( .A(n30506), .ZN(p_wishbone_bd_ram_n22619) );
  INV_X1 U34978 ( .A(n60975), .ZN(n30508) );
  INV_X1 U34979 ( .A(n30508), .ZN(p_wishbone_bd_ram_n22618) );
  INV_X1 U34980 ( .A(n60974), .ZN(n30510) );
  INV_X1 U34981 ( .A(n30510), .ZN(p_wishbone_bd_ram_n22617) );
  INV_X1 U34982 ( .A(n60973), .ZN(n30512) );
  INV_X1 U34983 ( .A(n30512), .ZN(p_wishbone_bd_ram_n22616) );
  INV_X1 U34984 ( .A(n60972), .ZN(n30514) );
  INV_X1 U34985 ( .A(n30514), .ZN(p_wishbone_bd_ram_n22615) );
  INV_X1 U34986 ( .A(n60971), .ZN(n30516) );
  INV_X1 U34987 ( .A(n30516), .ZN(p_wishbone_bd_ram_n22614) );
  INV_X1 U34988 ( .A(n60970), .ZN(n30518) );
  INV_X1 U34989 ( .A(n30518), .ZN(p_wishbone_bd_ram_n22613) );
  INV_X1 U34990 ( .A(n60969), .ZN(n30520) );
  INV_X1 U34991 ( .A(n30520), .ZN(p_wishbone_bd_ram_n22612) );
  INV_X1 U34992 ( .A(n60968), .ZN(n30522) );
  INV_X1 U34993 ( .A(n30522), .ZN(p_wishbone_bd_ram_n22611) );
  INV_X1 U34994 ( .A(n60967), .ZN(n30524) );
  INV_X1 U34995 ( .A(n30524), .ZN(p_wishbone_bd_ram_n22610) );
  INV_X1 U34996 ( .A(n60966), .ZN(n30526) );
  INV_X1 U34997 ( .A(n30526), .ZN(p_wishbone_bd_ram_n22609) );
  INV_X1 U34998 ( .A(n60965), .ZN(n30528) );
  INV_X1 U34999 ( .A(n30528), .ZN(p_wishbone_bd_ram_n22608) );
  INV_X1 U35000 ( .A(n60964), .ZN(n30530) );
  INV_X1 U35001 ( .A(n30530), .ZN(p_wishbone_bd_ram_n22607) );
  INV_X1 U35002 ( .A(n60963), .ZN(n30532) );
  INV_X1 U35003 ( .A(n30532), .ZN(p_wishbone_bd_ram_n22606) );
  INV_X1 U35004 ( .A(n60962), .ZN(n30534) );
  INV_X1 U35005 ( .A(n30534), .ZN(p_wishbone_bd_ram_n22605) );
  INV_X1 U35006 ( .A(n60961), .ZN(n30536) );
  INV_X1 U35007 ( .A(n30536), .ZN(p_wishbone_bd_ram_n22604) );
  INV_X1 U35008 ( .A(n60960), .ZN(n30538) );
  INV_X1 U35009 ( .A(n30538), .ZN(p_wishbone_bd_ram_n22603) );
  INV_X1 U35010 ( .A(n60959), .ZN(n30540) );
  INV_X1 U35011 ( .A(n30540), .ZN(p_wishbone_bd_ram_n22602) );
  INV_X1 U35012 ( .A(n60958), .ZN(n30542) );
  INV_X1 U35013 ( .A(n30542), .ZN(p_wishbone_bd_ram_n22601) );
  INV_X1 U35014 ( .A(n60957), .ZN(n30544) );
  INV_X1 U35015 ( .A(n30544), .ZN(p_wishbone_bd_ram_n22600) );
  INV_X1 U35016 ( .A(n60956), .ZN(n30546) );
  INV_X1 U35017 ( .A(n30546), .ZN(p_wishbone_bd_ram_n22599) );
  INV_X1 U35018 ( .A(n60955), .ZN(n30548) );
  INV_X1 U35019 ( .A(n30548), .ZN(p_wishbone_bd_ram_n22598) );
  INV_X1 U35020 ( .A(n60954), .ZN(n30550) );
  INV_X1 U35021 ( .A(n30550), .ZN(p_wishbone_bd_ram_n22597) );
  INV_X1 U35022 ( .A(n60953), .ZN(n30552) );
  INV_X1 U35023 ( .A(n30552), .ZN(p_wishbone_bd_ram_n22596) );
  INV_X1 U35024 ( .A(n60952), .ZN(n30554) );
  INV_X1 U35025 ( .A(n30554), .ZN(p_wishbone_bd_ram_n22595) );
  INV_X1 U35026 ( .A(n60951), .ZN(n30556) );
  INV_X1 U35027 ( .A(n30556), .ZN(p_wishbone_bd_ram_n22594) );
  INV_X1 U35028 ( .A(n60950), .ZN(n30558) );
  INV_X1 U35029 ( .A(n30558), .ZN(p_wishbone_bd_ram_n22593) );
  INV_X1 U35030 ( .A(n60949), .ZN(n30560) );
  INV_X1 U35031 ( .A(n30560), .ZN(p_wishbone_bd_ram_n22592) );
  INV_X1 U35032 ( .A(n60948), .ZN(n30562) );
  INV_X1 U35033 ( .A(n30562), .ZN(p_wishbone_bd_ram_n22591) );
  INV_X1 U35034 ( .A(n60947), .ZN(n30564) );
  INV_X1 U35035 ( .A(n30564), .ZN(p_wishbone_bd_ram_n22590) );
  INV_X1 U35036 ( .A(n60946), .ZN(n30566) );
  INV_X1 U35037 ( .A(n30566), .ZN(p_wishbone_bd_ram_n22589) );
  INV_X1 U35038 ( .A(n60945), .ZN(n30568) );
  INV_X1 U35039 ( .A(n30568), .ZN(p_wishbone_bd_ram_n22588) );
  INV_X1 U35040 ( .A(n60944), .ZN(n30570) );
  INV_X1 U35041 ( .A(n30570), .ZN(p_wishbone_bd_ram_n22587) );
  INV_X1 U35042 ( .A(n60943), .ZN(n30572) );
  INV_X1 U35043 ( .A(n30572), .ZN(p_wishbone_bd_ram_n22586) );
  INV_X1 U35044 ( .A(n60942), .ZN(n3